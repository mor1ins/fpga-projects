library ieee;
use ieee.std_logic_1164.all;
entity top is
    port
    (
        -- IN
        ------------------------------------------------------------------------------------------------------------------------------------------------------
        csi2_dphy_reset_n_i         : in std_logic; --         Asynchronous system reset (active low)
        csi2_dphy_reset_byte_fr_n_i : in std_logic; --         Active low reset. Resets the nets in the clk_byte_fr clock domain. The signal driving this
        --                                                              port must already be synchronized to the clk_byte_fr. 
        csi2_dphy_reset_byte_n_i : in std_logic; --            Active low reset. Resets the logic clocked by the clk_byte_o.
        csi2_dphy_reset_lp_n_i   : in std_logic; --            Active low reset. This resets the nets in the clk_lp_hs_ctrl clock domain. The signal
        --                                                              driving this port must already be synchronized to the clk_lp_hs_ctrl. No need to drive
        --                                                              this reset if the Rx clock mode is HS_ONLY.

        csi2_dphy_clk_byte_fr_i : in std_logic; --             Continuously running byte clock. This should be div8 (in gear16) or div4 (in gear8) of the
        --                                                              input D-PHY clock. This also clocks the logic that detects the Rx D-PHY data lane
        --                                                              transitions (lp_hs_ctrl_d0-3 modules). This is also used by the word_align, lane_align
        --                                                              and capture_control modules. Payload output is also in this clock domain
        csi2_dphy_clk_lp_ctrl_i : in std_logic; --             Clocks the logic that detects the Low Power states of the D-PHY clock lane. The period of
        --                                                              this clock should be smaller than the tLPX, with enough setup and hold time, to properly sample
        --                                                              the Low Power state transitions. No need to drive this reset if the Rx clock mode is HS_ONLY.

        csi2_dphy_pd_dphy_i  : in std_logic; --                Active high. Power Down control signal. Applicable only for Hard D-PHY implementation.
        csi2_dphy_pll_lock_i : in std_logic; --                PLL lock indicator, if a PLL is used to generate a free-running byte clock. Set this to 1 if a
        --                                                              PLL is not used. Active high.
        ------------------------------------------------------------------------------------------------------------------------------------------------------

        -- OUT
        ------------------------------------------------------------------------------------------------------------------------------------------------------
        csi2_dphy_bd0_o : out std_logic_vector(7 downto 0); --      Byte Data directly from lane 0. This is 8-bit wide for gear 8, 16 bits for gear 16

        csi2_dphy_lp_hs_state_clk_o : out std_logic_vector(1 downto 0); --     2-bit state encoding of the D-PHY clock controller
        csi2_dphy_lp_hs_state_d_o   : out std_logic_vector(1 downto 0); --     2-bit state encoding of the D-PHY data lane 0 controller

        csi2_dphy_clk_byte_hs_o : out std_logic; --         Generated byte clock from the D-PHY module based on the input D-PHY clock lane,
        --                                                              active only when the clock lanes are in high-speed mode. This clock is the same as the
        --                                                              clk_byte_o when the submodule is in HS_ONLY mode and D-PHY implementation is Soft DPHY.
        --                                                              This may be connected to the clk_byte_fr_i when the RX Clock Mode is HS_ONLY.
        csi2_dphy_clk_byte_o : out std_logic; --            Generated byte clock from the D-PHY module based on the input D-PHY clock lane, used
        --                                                              to latch the internal parallel byte data from dphy_rx_wrap. This is div4 or div8 of the
        --                                                              D-PHY clock lane frequency. This is only active when the data lanes are in high-speed mode

        csi2_dphy_capture_en_o : out std_logic; --          Indicates valid byte data in bd0/1/2/3_o.
        csi2_dphy_cd_d0_o      : out std_logic; --          Contention detection indicator. Active high.

        csi2_dphy_hs_d_en_o : out std_logic; --             Active-high high-speed mode enable for data lane d0. For Hard D-PHY IP, this signal is
        --                                                              also used for HS mode enable for the other data lanes.
        csi2_dphy_hs_sync_o : out std_logic; --             This indicates the successful detection of the synchronization code ‘B8 in the data lanes.
        --                                                              This signal asserts from the start of synchronization pattern ‘B8 up to the last data
        --                                                              captured before detecting LP-11 state (of any lane, if Soft D-PHY; of data lane0 for Hard
        --                                                              D-PHY). Active high.
        csi2_dphy_lp_d0_rx_n_o : out std_logic; --          Low-power values of data lane 0 true and differential lines, respectively.
        csi2_dphy_lp_d0_rx_p_o : out std_logic;

        csi2_dphy_term_clk_en_o : out std_logic; --          Active-high enable signal for the line termination of the D-PHY clock lane. This is
        --                                                              asserted on detection of transition from LP-11 to LP-01 of the clock lane, and deasserts
        --                                                              upon detection of LP-11 after a high-speed mode.
        ------------------------------------------------------------------------------------------------------------------------------------------------------

        -- INOUT
        ------------------------------------------------------------------------------------------------------------------------------------------------------
        csi2_dphy_clk_n_i : inout std_logic; --             MIPI D-PHY clock lane
        csi2_dphy_clk_p_i : inout std_logic; --             MIPI D-PHY clock lane

        csi2_dphy_d0_n_i : inout std_logic; --              MIPI D-PHY data lane 0. Available only for MIPI CSI-2 configuration.
        csi2_dphy_d0_p_i : inout std_logic  --               MIPI D-PHY data lane 0. Available only for MIPI CSI-2 configuration.
        ------------------------------------------------------------------------------------------------------------------------------------------------------
    );
end entity top; -- sbp_module=true 

architecture rtl of top is
    component csi2_dphy is
        port
        (
            bd0_o             : out std_logic_vector(7 downto 0);
            lp_hs_state_clk_o : out std_logic_vector(1 downto 0);
            lp_hs_state_d_o   : out std_logic_vector(1 downto 0);
            capture_en_o      : out std_logic;
            cd_d0_o           : out std_logic;
            clk_byte_fr_i     : in std_logic;
            clk_byte_hs_o     : out std_logic;
            clk_byte_o        : out std_logic;
            clk_lp_ctrl_i     : in std_logic;
            clk_n_i           : inout std_logic;
            clk_p_i           : inout std_logic;
            d0_n_i            : inout std_logic;
            d0_p_i            : inout std_logic;
            hs_d_en_o         : out std_logic;
            hs_sync_o         : out std_logic;
            lp_d0_rx_n_o      : out std_logic;
            lp_d0_rx_p_o      : out std_logic;
            pll_lock_i        : in std_logic;
            reset_byte_fr_n_i : in std_logic;
            reset_byte_n_i    : in std_logic;
            reset_lp_n_i      : in std_logic;
            reset_n_i         : in std_logic;
            term_clk_en_o     : out std_logic
        );

    end component csi2_dphy; -- not_need_bbox=true 

begin
    csi2_dphy_inst : component csi2_dphy port map
    (
        bd0_o(7)      => csi2_dphy_bd0_o(7),
        bd0_o(6) => csi2_dphy_bd0_o(6), bd0_o(5) => csi2_dphy_bd0_o(5), bd0_o(4) => csi2_dphy_bd0_o(4),
        bd0_o(3) => csi2_dphy_bd0_o(3), bd0_o(2) => csi2_dphy_bd0_o(2), bd0_o(1) => csi2_dphy_bd0_o(1),
        bd0_o(0) => csi2_dphy_bd0_o(0), lp_hs_state_clk_o(1) => csi2_dphy_lp_hs_state_clk_o(1),
        lp_hs_state_clk_o(0) => csi2_dphy_lp_hs_state_clk_o(0), lp_hs_state_d_o(1) => csi2_dphy_lp_hs_state_d_o(1),
        lp_hs_state_d_o(0) => csi2_dphy_lp_hs_state_d_o(0), capture_en_o => csi2_dphy_capture_en_o,
        cd_d0_o => csi2_dphy_cd_d0_o, clk_byte_fr_i => csi2_dphy_clk_byte_fr_i,
        clk_byte_hs_o => csi2_dphy_clk_byte_hs_o, clk_byte_o => csi2_dphy_clk_byte_o,
        clk_lp_ctrl_i => csi2_dphy_clk_lp_ctrl_i, clk_n_i => csi2_dphy_clk_n_i,
        clk_p_i => csi2_dphy_clk_p_i, d0_n_i => csi2_dphy_d0_n_i, d0_p_i => csi2_dphy_d0_p_i,
        hs_d_en_o => csi2_dphy_hs_d_en_o, hs_sync_o => csi2_dphy_hs_sync_o,
        lp_d0_rx_n_o => csi2_dphy_lp_d0_rx_n_o, lp_d0_rx_p_o => csi2_dphy_lp_d0_rx_p_o, pll_lock_i => csi2_dphy_pll_lock_i,
        reset_byte_fr_n_i => csi2_dphy_reset_byte_fr_n_i, reset_byte_n_i => csi2_dphy_reset_byte_n_i,
        reset_lp_n_i => csi2_dphy_reset_lp_n_i, reset_n_i => csi2_dphy_reset_n_i,
        term_clk_en_o => csi2_dphy_term_clk_en_o);

end architecture rtl; -- sbp_module=true 