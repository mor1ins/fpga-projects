module gamma_correction (
     r_in,
     g_in,
     b_in,
	 
     r_out,
     g_out,
     b_out
);


input [11:0] r_in, g_in, b_in;
output [11:0] r_out, g_out, b_out;




endmodule  