// =========================================================================
// Filename: byte2pixel_tb.v
// Copyright(c) 2019 Lattice Semiconductor Corporation. All rights reserved.
// =========================================================================

////////////////////////////////////////////////////////
/// � Intermotion Technology
/// � B2P Changes
/// � Date MAY 2, 2019
/// � Arman Arshakyan
/// � Some directives are changed to parameters.
/// � Changed/updated some signals/parameters names.
/// � Changed/updated some structural solutions.
/// � Added solution to automatically compare data files "expected_data.log" vs "received_data.log" and "expected_sync_data.log" vs "received_sync_data.log".  
//////////////////////////////////////////////////////////////////////////////////

#include <orcapp_head>
`timescale 1 ps / 1 ps

`include "tb_defs.v"
`include "byte_driver.v"
`include "pixel_monitor.v"

`ifndef NUM_FRAMES
  `define NUM_FRAMES 1
`endif
`ifndef NUM_LINES 
  `define NUM_LINES 1
`endif
`ifndef NUM_BYTES
  `define NUM_BYTES 180
`endif
`ifndef HFP_PAYLOAD
  `define HFP_PAYLOAD 110
`endif
`ifndef HSA_PAYLOAD
  `define HSA_PAYLOAD 40
`endif
`ifndef HBP_PAYLOAD
  `define HBP_PAYLOAD 220
`endif
`ifndef VFP_LINES
  `define VFP_LINES 5
`endif
`ifndef VSA_LINES
  `define VSA_LINES 5
`endif
`ifndef VBP_LINES
  `define VBP_LINES 20
`endif

module byte2pixel_tb;
`include "dut_params.v"
`include "test_dsi_reset.v" 
`include "test_csi2_reset.v" 
     
   PUR PUR_INST(.PUR(1'b1));
   GSR GSR_INST(.GSR(1'b1));

localparam RGB666          = 6'h1E;
localparam RGB666_LOOSE    = 6'h2E;
localparam RAW8            = 6'h2A;
localparam RAW10           = 6'h2B;
localparam RAW12           = 6'h2C;
localparam YUV420_8        = 6'h18;
localparam YUV420_8_CSPS   = 6'h1C;
localparam LEGACY_YUV420_8 = 8'h1A;
localparam YUV422_8        = 8'h1E;
localparam YUV420_10       = 8'h19;
localparam YUV420_10_CSPS  = 8'h1D;
localparam YUV422_10       = 8'h1F;
localparam RGB888          = (RX_TYPE=="DSI") ? 6'h3E : 6'h24;
 
localparam DT =     (DATA_TYPE == "RGB888")          ? RGB888 :
                    (DATA_TYPE == "RGB666")          ? RGB666 :
                    (DATA_TYPE == "RGB666_LOOSE")    ? RGB666_LOOSE :
                    (DATA_TYPE == "RAW8")            ? RAW8 :
                    (DATA_TYPE == "RAW10")           ? RAW10 :
                    (DATA_TYPE == "RAW12")           ? RAW12 :
                    (DATA_TYPE == "YUV420_8")        ? YUV420_8 :
                    (DATA_TYPE == "YUV420_8_CSPS")   ? YUV420_8_CSPS :
                    (DATA_TYPE == "LEGACY_YUV420_8") ? LEGACY_YUV420_8 :
                    (DATA_TYPE == "YUV422_8")        ? YUV422_8 :
                    (DATA_TYPE == "YUV420_10")       ? YUV420_10 :
                    (DATA_TYPE == "YUV420_10_CSPS")  ? YUV420_10_CSPS :
                    (DATA_TYPE == "YUV422_10")       ? YUV422_10 : RGB888;

localparam BWIDTH = (DATA_TYPE == "RGB888")          ? 24 :
                    (DATA_TYPE == "RGB666")          ? 18 :
                    (DATA_TYPE == "RGB666_LOOSE")    ? 18 :
                    (DATA_TYPE == "RAW8")            ?  8 :
                    (DATA_TYPE == "RAW10")           ? 10 :
                    (DATA_TYPE == "RAW12")           ? 12 :
                    (DATA_TYPE == "YUV420_8")        ?  8 :
                    (DATA_TYPE == "YUV420_8_CSPS")   ?  8 :
                    (DATA_TYPE == "LEGACY_YUV420_8") ?  8 :
                    (DATA_TYPE == "YUV422_8")        ?  8 :
                    (DATA_TYPE == "YUV420_10")       ? 10 :
                    (DATA_TYPE == "YUV420_10_CSPS")  ? 10 :
                    (DATA_TYPE == "YUV422_10")       ? 10 : 24;

localparam LOOSE_CNT      = PD_BUS_WIDTH/BWIDTH;
`ifdef SIP_PCLK
localparam PIXCLK_PERIOD  = `SIP_PCLK/2;
`else
localparam PIXCLK_PERIOD  = (DATA_TYPE == "RGB666_LOOSE") ? `SIP_BCLK*24*LOOSE_CNT*NUM_TX_CH/(2*NUM_RX_LANE*RX_GEAR) :
                                                            `SIP_BCLK*PD_BUS_WIDTH*NUM_TX_CH/(2*NUM_RX_LANE*RX_GEAR) ;
`endif

parameter BYTECLK_PERIOD  = `SIP_BCLK/2;
//parameter NUM_BYTES       = `NUM_BYTES;
parameter NUM_BYTES       = PD_BUS_WIDTH * 48;
parameter NUM_LINES       = `NUM_LINES;
parameter NUM_FRAMES      = `NUM_FRAMES;
parameter PIXEL_COUNT     = PD_BUS_WIDTH*NUM_TX_CH/BWIDTH;

`ifdef SP2_LP_SIMULTANEOUS
parameter SP2_LP_ENABLE   = 1;
parameter SP_LP2_ENABLE   = 0;
`elsif SP_LP2_SIMULTANEOUS
parameter SP_LP2_ENABLE   = 1;
parameter SP2_LP_ENABLE   = 0;
`else                         
parameter SP2_LP_ENABLE   = 0;
parameter SP_LP2_ENABLE   = 0;
`endif

reg                                 reset_byte_n_i;
reg                                 reset_pixel_n_i;
reg                                 clk_byte_i;
reg                                 clk_pixel_i;
wire [5:0]                          dt_i;
wire [5:0]                          dt2_i;
wire                                sp_en_i;
wire                                sp2_en_i;
wire                                lp_av_en_i;
wire                                lp2_av_en_i;
wire [(RX_GEAR*NUM_RX_LANE)-1:0]    payload_i ;
wire                                payload_en_i;
wire [15:0]                         wc_i;
wire [15:0]                         wc2_i;
wire [(PD_BUS_WIDTH*NUM_TX_CH)-1:0] pd_o;
wire [1:0]p_odd_o;
wire hsync_o, vsync_o, fv_o, lv_o, de_o;
wire hsync_w, vsync_w, fv_w, lv_w, de_w;
wire [3:0]                        write_cycle_o;  
wire                              mem_we_o;       
wire                              mem_re_o;       
wire [1:0]                        read_cycle_o;   
wire [2:0]                        mem_radr_o;     

reg                  start_video      = 0;
reg                  enable_write_log = 1;
reg [4:0]            wait_cycles;
reg                  error_flag;
reg                  p_odd_error_flag;
reg [PD_BUS_WIDTH:0] expected_data;
reg [PD_BUS_WIDTH:0] received_data;
reg [5*8-1:0]        expected_sync;
reg [5*8-1:0]        received_sync;
integer              comp_pixel_num;
integer              pixel_count_error;
integer              pixel_mismatch_counter;
integer              comp_sync_num;
integer              sync_count_error;
integer              sync_mismatch_counter;
integer              sync_in_file;
integer              sync_out_file;
integer              expected_file; // file handler
integer              received_file; // file handler
integer              scan_in_file; // file handler
integer              scan_out_file; // file handler

//BYTE RESET LOGIC
    initial begin
        reset_byte_n_i  = 1;
        reset_pixel_n_i = 1;
        repeat(3) @(posedge clk_byte_i)
        reset_byte_n_i  = 0;
        reset_pixel_n_i = 0;
        repeat(4) @(posedge clk_pixel_i)
        reset_byte_n_i  = 1;
        reset_pixel_n_i = 1;
    end

    initial begin
        clk_pixel_i= 1;
        forever begin
            #PIXCLK_PERIOD clk_pixel_i= ~clk_pixel_i;
        end
    end

    initial begin
        clk_byte_i = 1;
        forever begin
            #BYTECLK_PERIOD clk_byte_i = ~clk_byte_i;
        end
    end
//--------------------------------------------------------------------------------------------------

// USERNAME byte2pixel_dut(
//                    .reset_byte_n_i      (reset_byte_n_i),
//                    .clk_byte_i          (clk_byte_i),
//                    .sp_en_i             (sp_en_i),       // Short Packet Enable
//                    .sp2_en_i            (sp2_en_i),      // Short Packet Enable #2
//                    .dt_i                (dt_i),       // Data Type
//                    .dt2_i               (dt2_i),      // Data Type #2
//                    .lp_av_en_i          (lp_av_en_i),        // Long Packet of Active Video Enable
//                    .lp2_av_en_i         (lp2_av_en_i),       // Long Packet of Active Video Enable #2
//                    .payload_en_i        (payload_en_i),      // paload enable
//                    .payload_i           (payload_i),         // payload_i
//                    .wc_i                (wc_i),        // payload_i byte count
//                    .wc2_i               (wc2_i),       // payload_i byte count #2
//                    .reset_pixel_n_i     (reset_pixel_n_i),
//                    .clk_pixel_i         (clk_pixel_i),   
//                    //outputs
//                    .vsync_o             (vsync_o),         // Vsync in clk_pixel domain
//                    .hsync_o             (hsync_o),         // Hsync in clk_pixel domain
//                    .fv_o                (fv_o),            // Frame Valid in clk_pixel domain
//                    .lv_o                (lv_o),            // Line Valid in clk_pixel_i domain
//                    .de_o                (de_o),            // picture data enable
//                    .pd_o                (pd_o),            // picture data
//                                                            
//                    .p_odd_o             (p_odd_o),         // odd pixel indicator
//                    .write_cycle_o       ( ),               // payload_i Write Cycle (for debug)
//                    .mem_we_o            ( ),               // payload_i Write Enable (for debug)
//                    .mem_re_o            ( ),               // payload_i Read Enable (for debug)
//                    .read_cycle_o        ( ),               // pixel data Read Cycle (for debug)
//                    .mem_radr_o          ( )                // pixel data Read Address (for debug)
//                   );
//--------------------------------------------------------------------------------------------------
`include "dut_inst.v"

     byte_driver #(
                   .DATA_TYPE            (DT),
                   .RX_TYPE              (RX_TYPE),
                   .DSI_MODE             (DSI_MODE),
                   .GEAR                 (RX_GEAR),
                   .RX_CH                (NUM_RX_LANE),
                   .PD_BUS_WIDTH         (PD_BUS_WIDTH),
                   .NUM_TX_CH            (NUM_TX_CH),
                   .NUM_BYTES            (NUM_BYTES),
                   .NUM_LINES            (NUM_LINES),
                   .SP_LP2_ENABLE        (SP_LP2_ENABLE),
                   .SP2_LP_ENABLE        (SP2_LP_ENABLE)
                  )
    u_data_driver (
                   .enable_write_log     (enable_write_log),
                   .hsync_o              (hsync_o),
                   .clk                  (clk_byte_i),
                   .reset                (~reset_byte_n_i),
                   .vid_cntl_tgen_active (start_video),
                   .sp_o                 (sp_en_i),
                   .lp_o                 (lp_av_en_i),
                   .dt_o                 (dt_i),
                   .wc_o                 (wc_i),
                   .sp2_o                (sp2_en_i),
                   .lp2_o                (lp2_av_en_i),
                   .dt2_o                (dt2_i),
                   .wc2_o                (wc2_i),
                   .payload_en           (payload_en_i),
                   .byte_data            (payload_i)
                  );
//--------------------------------------------------------------------------------------------------

assign vsync_w      = (CTRL_POL == "POSITIVE") ? vsync_o : ~vsync_o;
assign hsync_w      = (CTRL_POL == "POSITIVE") ? hsync_o : ~hsync_o;
assign de_w         = (CTRL_POL == "POSITIVE") ? de_o    : ~de_o;
assign fv_w         = (CTRL_POL == "POSITIVE") ? fv_o    : ~fv_o;
assign lv_w         = (CTRL_POL == "POSITIVE") ? lv_o    : ~lv_o;

    pixel_monitor #(
                   .RX_TYPE         (RX_TYPE),
                   .PD_BUS_WIDTH    (PD_BUS_WIDTH),
                   .PIXEL_COUNT     (PIXEL_COUNT),
                   .TX_CH           (NUM_TX_CH)
                   )
    u_pixel_monitor (
                   .enable_write_log (enable_write_log),
                   .clk              (clk_pixel_i),
                   .reset            (~reset_pixel_n_i),
                   .vsync            (vsync_w),
                   .hsync            (hsync_w),
                   .de_o             (de_w),
                   .frame_valid      (fv_w),
                   .line_valid       (lv_w),
                   .pixel_data       (pd_o)
                  );

 // reset tests
`ifdef DSI_RESET_DE
    initial begin
        dsi_reset_de; //call the task
    end
`elsif DSI_RESET_HSYNC
    initial begin
        dsi_reset_hsync; //call the task
    end
`elsif DSI_RESET_VSYNC
    initial begin
        dsi_reset_vsync; //call the task
    end
`elsif DSI_RESET_DE_NEG
    initial begin
        dsi_reset_de_neg; //call the task
    end
`elsif DSI_RESET_HSYNC_NEG
    initial begin
        dsi_reset_hsync_neg; //call the task
    end
`elsif DSI_RESET_VSYNC_NEG
    initial begin
        dsi_reset_vsync_neg; //call the task
    end
`elsif CSI2_RESET_FV
    initial begin
        csi_reset_fv;
    end
`elsif CSI2_RESET_LV
    initial begin
        csi_reset_lv;
    end
`else

// clean off the content of existing files if any
    initial begin
        if(enable_write_log == 1) begin
            expected_file = $fopen("expected_data.log","w");
            $fclose(expected_file);

            received_file = $fopen("received_data.log","w");
            $fclose(received_file);
            
            if (RX_TYPE == "DSI") begin
                sync_in_file = $fopen("expected_sync_data.log","w");
                $fclose(sync_in_file);
            
                sync_out_file = $fopen("received_sync_data.log","w");
                $fclose(sync_out_file);
            end
        end
    end
    
    initial begin
        `define NULL 0
        start_video = 1;
        error_flag = 0;
        comp_pixel_num = 0;
        pixel_count_error = 0;
        pixel_mismatch_counter = 0;
        comp_sync_num = 0;
        sync_mismatch_counter = 0;

        @(posedge reset_pixel_n_i) 
        $display ("******************************");
        $display (">>>>> TRANSMITTING DATA <<<<< ");
        if (RX_TYPE == "DSI") 
            repeat(NUM_FRAMES+1) @(negedge vsync_w);
        else //(RX_TYPE == "CSI2") 
            repeat(NUM_FRAMES) @(negedge fv_w);
        #100; 
        $display ("-----------------------------");
        $display (">>>>> TRANSMIT DONE !!! <<<<<");
        $display ("*****************************");

        if(enable_write_log == 1) begin
// Data comparing
            expected_file = $fopen("expected_data.log", "r");
            received_file = $fopen("received_data.log", "r");
            if (expected_file == `NULL) begin
                $display (">>>>> E R R O R : expected_data.log file handle was NULL");
                $finish;
            end
            if (received_file == `NULL) begin
                $display (">>>>> E R R O R : received_data.log file handle was NULL");
                $finish;
            end
            $display ("----------------------------------------------------------------------------------------------------------");
            $display (">>>>> I N F O   : Expected and Received Pixel Data are saved in expected_data.log and received_data.log!!!");
            $display ("----------------------------------------------------------------------------------------------------------");
            
            $display ("---------------------------------------------------------------------");
            $display (">>>>> I N F O   : PIXEL DATA COMPARISON -> EXPECTED vs RECEIVED <<<<<");
            $display ("---------------------------------------------------------------------");
            if (u_data_driver.expected_pixel_counter != u_pixel_monitor.received_pixel_counter) begin
            error_flag = 1;
            end
            while (!$feof(expected_file) && !$feof(received_file)) begin
                scan_in_file  = $fscanf(expected_file, "%h\n", expected_data);
                scan_out_file = $fscanf(received_file, "%h\n", received_data);
                comp_pixel_num = comp_pixel_num +1;
                if (expected_data !== received_data) begin
                    $display (">>>>> E R R O R : Expected and Received pixel data mismatch. Line %0d", comp_pixel_num);
                    $display ("       Expected:  %h", expected_data);
                    $display ("       Received:  %h", received_data);
                    error_flag = 1;
                    pixel_mismatch_counter = pixel_mismatch_counter + 1;
                end
            end
        
            if (pixel_mismatch_counter > 0) begin
//                $display("**** I N F O : Actual Pixel Count is %0d", actual_pixel_counter);
//                $display("**** I N F O : Expected Pixel Count is %0d", exp_pixel_count);
                $display (">>>>> I N F O   : Pixels Mismatch Count=%0d", pixel_mismatch_counter);
                $display ("-------------------------------------------");
                error_flag = 1;
            end
        
            if ($feof(expected_file) && $feof(received_file)) begin
                $display (">>>>> I N F O   : Expected and Rceived pixel counts are equal");
            end
            else begin 
                $display (">>>>> E R R O R : Expected and Rceived pixel counts are not equal");
                pixel_count_error = 1;
                error_flag = 1;
            end   
        
            $display (">>>>> I N F O   : Expected Pixel count=%0d", u_data_driver.expected_pixel_counter);
            $display (">>>>> I N F O   : Received Pixel count=%0d", u_pixel_monitor.received_pixel_counter);
            $display ("---------------------------------------------------------------");
            $display (">>>>> I N F O   : NUM_FRAMES=%0d, NUM_LINES=%0d, Word Count=%0d", NUM_FRAMES, NUM_LINES, NUM_BYTES);
            $display ("---------------------------------------------------------------");

// hsync/vsync data comparing
            if (RX_TYPE == "DSI") begin
                sync_in_file  = $fopen("expected_sync_data.log", "r");
                sync_out_file = $fopen("received_sync_data.log", "r");
                if (sync_in_file == `NULL) begin
                    $display (">>>>> E R R O R : expected_sync_data.log file handle was NULL");
                end
                if (sync_out_file == `NULL) begin
                    $display (">>>>> E R R O R : received_sync_data.log file handle was NULL");
                end
                $display ("---------------------------------------------------------------------------------------------------------------------------");
                $display (">>>>> I N F O   : Expected and Received HSYNC/VSYNC Datas are saved in expected_sync_data.log and received_sync_data.log!!!");
                $display ("---------------------------------------------------------------------------------------------------------------------------");
            
                while (!$feof(sync_in_file) && !$feof(sync_out_file)) begin
                    scan_in_file  = $fscanf(sync_in_file, "%s\n", expected_sync);
                    scan_out_file = $fscanf(sync_out_file, "%s\n", received_sync);
                    comp_sync_num = comp_sync_num + 1;
                    if (expected_sync !== received_sync) begin
                        $display (">>>>> E R R O R : Expected and Received hsync/vsync data mismatch. Line %0d", comp_sync_num);
                        $display ("       Expected:  %s", expected_sync);
                        $display ("       Received:  %s", received_sync);
                        error_flag = 1;
                        sync_mismatch_counter = sync_mismatch_counter + 1;
                    end
                end
                if (sync_mismatch_counter > 0) begin
                    $display (">>>>> I N F O   : hsync/vsync Mismatch Count=%0d", sync_mismatch_counter);
                    $display ("------------------------------------------------");
                    error_flag = 1;
                end
                if ($feof(sync_in_file) && $feof(sync_out_file)) begin
                    $display (">>>>> I N F O   : Expected and Rceived hsinc/vsync counts are equal");
                    $display (">>>>> I N F O   : hsinc/vsync count=%0d", comp_sync_num);
                    $display ("-------------------------------------------------------------------");
                end
                else begin 
                    $display (">>>>> E R R O R : Expected and Rceived hsinc/vsync counts are not equal");
                    $display ("-----------------------------------------------------------------------");
                    sync_count_error = 1;
                    error_flag = 1;
                end   
            end
            
            if (error_flag == 1) begin
                if (p_odd_error_flag == 1) begin
                    $display (">>>>> E R R O R : p_odd_o signal is x/z");
                    $display ("---------------------------------------");
                end 
                $display ("********** T E S T     F A I L E D **********");
                $display ("---------------------------------------------");
            end
            else begin
                $display ("********** SIMULATION PASSED **********");
                $display ("--------------------------------------");
            end
            $finish;
        end
    end
`endif

    initial begin
        if (RX_TYPE == "DSI") 
            dsi_default_val_check;
        else //(RX_TYPE == "CSI2")
            csi_default_val_check;
    end

generate
  if (RX_TYPE=="DSI") begin
    initial begin
        forever begin
            @(posedge reset_pixel_n_i);
            #1;
            if( |p_odd_o === 1'bx || |p_odd_o === 1'bz) begin
//                $display (">>>>> E R R O R : p_odd_o signal is x/z");
//                $display ("---------------------------------------");
                p_odd_error_flag = 1;
                error_flag = 1;
                //#1000 $finish;
            end
        end
    end
  end
endgenerate

endmodule
