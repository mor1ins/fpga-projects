`define DEVICE_ECP5U   
`timescale 1ns/100ps
module colorspace (
               clk,
               din0,
               din1,
               din2,
               dout0,
               dout1,
               dout2,
               rstn
        );
   input                         rstn ;
   input                         clk ;
   input  [12-1:0]  din0;
   input  [12-1:0]  din1;
   input  [12-1:0]  din2;
   output [12-1:0] dout0; 
   output [12-1:0] dout1; 
   output [12-1:0] dout2; 
 csc_core_colorspace #(.CORETYPE          (0),
              .CWIDTH            (9),
              .CPOINTS           (7),
              .DINWIDTH          (12),
              .DINSIGN           ("Unsigned"),
              .DOUTWIDTH         (12),
              .DOUTPOINTS        (0),
              .DOUTSIGN          ("Unsigned"),
              .LSBMETHOD         ("Rounding up"),
              .MSBMETHOD         ("Saturation"),
              .INREG             ("Enable"),
              .IOVALID           (0),
              .INSERIAL          ("Parallel"),
              .DSPBLKMULT        ("Disable"),
              .TAGSWIDTH         (1),
              .LATENCY           (9),
              .CV_MH             (9'h080), 
              .CV_MI             (9'h000), 
              .CV_MJ             (9'h000), 
              .CV_MK             (21'h000000), 
              .CV_NH             (9'h000), 
              .CV_NI             (9'h080), 
              .CV_NJ             (9'h000), 
              .CV_NK             (21'h000000), 
              .CV_PH             (9'h000), 
              .CV_PI             (9'h000), 
              .CV_PJ             (9'h080), 
              .CV_PK             (21'h000000), 
              .DEVICE            ("ECP5U"),
              .OPTIMIZE          (0))
u1_core (
            .ce                  (1'b1          ),
            .sr                  (1'b0          ),
            .clk                 (clk           ),
            .inpvalid            (1'b1          ),
            .outvalid            (              ),
            .din0                (din0          ),
            .din1                (din1          ),
            .din2                (din2          ),
            .dout0               (dout0         ),
            .dout1               (dout1         ),
            .dout2               (dout2         ),
            .tags_in             (              ),
            .tags_out            (              ),
            .rstn                (rstn          )
         );
endmodule
// obf_with_line.v generated by Lattice IP Model Creator version 1
// created on Tue Feb 24 14:02:19 PST 2015
// Copyright(c) 2007 Lattice Semiconductor Corporation. All rights reserved
// obfuscator_exe version 1.mar0807
// top
module csc_core_colorspace (
               
               clk,              
               rstn,             
               ce,               
               sr,               
               inpvalid,         
               din0,                
               din1,             
               din2,             
               tags_in,          
               tags_out,         
               
               outvalid,         
               dout2,            
               dout1,            
               dout0             
               )
              `ifdef DEVICE_EC
               
              `else
               `ifdef DEVICE_ECP
                  
               `else
                  `ifdef DEVICE_ECP2
                     
                  `else
                     `ifdef DEVICE_ECP2M
                        
                     `else
                        `ifdef DEVICE_XP
                           
                        `else
                           `ifdef DEVICE_XP2
                              
                           `else
                              `ifdef DEVICE_SC
                                 
                              `else
                                 `ifdef DEVICE_SCM
                                    
                                 `else
                                    `ifdef DEVICE_ECP3
                                       
                                    `else
                                       `ifdef DEVICE_XO2
                                          
                                       `else
                                          `ifdef DEVICE_ECP5U
                                             
                                          `else
                                             `ifdef DEVICE_ECP5UM
                                                
                                             `else
                                                
                                             `endif
                                          `endif
                                       `endif
                                    `endif
                                 `endif
                              `endif
                           `endif
                        `endif
                     `endif
                  `endif
               `endif
            `endif
             
             ;
parameter   CORETYPE             =  0;
parameter   CWIDTH               =  8;
parameter   CPOINTS              =  0;
parameter   DINWIDTH             =  8;
parameter   DINSIGN              = "Signed";
parameter   DOUTWIDTH            =  8;
parameter   DOUTPOINTS           =  0;
parameter   DOUTSIGN             = "Signed";
parameter   LSBMETHOD            = "Rounding";
parameter   MSBMETHOD            = "Saturation";
parameter   INREG                = "Enbale";
parameter   INSERIAL             = "Serial";
parameter   KEEPBLANK            =  0;
parameter   DSPBLKMULT           = "Enable";
parameter   TAGSWIDTH            =  1;
parameter   IOVALID              =  1;
parameter   LATENCY              =  1;
parameter   CV_MH                =  0;
parameter   CV_MI                =  0;
parameter   CV_MJ                =  0;
parameter   CV_MK                =  0;
parameter   CV_NH                =  0;
parameter   CV_NI                =  0;
parameter   CV_NJ                =  0;
parameter   CV_NK                =  0;
parameter   CV_PH                =  0;
parameter   CV_PI                =  0;
parameter   CV_PJ                =  0;
parameter   CV_PK                =  0;
parameter   DEVICE               = "ECP2";
parameter   OPTIMIZE             =  0;
localparam ym3b97e          = DINWIDTH + CWIDTH;
localparam vk2fc20        = ym3b97e + 1;
localparam gof081f        = vk2fc20 + 1;
localparam je207ce               = rv3e73(LATENCY-1);
input                                  clk;
input                                  rstn;
input                                  ce;
input                                  sr;
input                                  inpvalid;
input  [DINWIDTH-1:0]                  din0;
input  [DINWIDTH-1:0]                  din1;
input  [DINWIDTH-1:0]                  din2;
input  [TAGSWIDTH-1:0]                 tags_in;
output                                 outvalid;
output [DOUTWIDTH-1:0]                 dout0;
output [DOUTWIDTH-1:0]                 dout1;
output [DOUTWIDTH-1:0]                 dout2;
output [TAGSWIDTH-1:0]                 tags_out;
wire   [gof081f-1:0]            cz51c7a;
wire   [gof081f-1:0]            th71ea7;
wire   [gof081f-1:0]            kd7a9fd;
wire   [DINWIDTH-1:0]                  pua7f60;
wire   [DINWIDTH-1:0]                  offd81a;
wire   [DINWIDTH-1:0]                  gb606af;
wire   [DINWIDTH-1:0]                  aa1abef;
wire   [DINWIDTH-1:0]                  rvafbca;
wire                                   ea7de57;
wire                                   meef2b9;
wire   [DINWIDTH-1:0]                  dmcae42;
wire   [DINWIDTH-1:0]                  gqb9092;
wire   [DINWIDTH-1:0]                  ne42486;
wire                                   gd12433;
wire                                   ec9219c;
wire   [DOUTWIDTH-1:0]                 hq86704;
wire   [DOUTWIDTH-1:0]                 ba9c11c;
wire   [DOUTWIDTH-1:0]                 ba4718;
wire   [TAGSWIDTH-1:0]                 zz1c615;
reg                                    lde30af;
reg                                    cb1857e;
wire   [DOUTWIDTH-1:0]                 uk15fae;
wire   [DOUTWIDTH-1:0]                 rt7eb87;
wire   [DOUTWIDTH-1:0]                 qvae1f1;
reg    [DOUTWIDTH-1:0]                 gq87c65;
reg    [DOUTWIDTH-1:0]                 byf1941;
reg    [DOUTWIDTH-1:0]                 uv6505b;
reg    [TAGSWIDTH-1:0]                 ip416ef;
reg ngb77c;
reg kd5bbe3;
reg vvddf1d;
reg [DINWIDTH - 1 : 0] jc7c771;
reg [DINWIDTH - 1 : 0] oh1dc57;
reg [DINWIDTH - 1 : 0] jp715e2;
reg [TAGSWIDTH - 1 : 0] jc578b4;
reg [gof081f - 1 : 0] ale2d18;
reg [gof081f - 1 : 0] qvb462f;
reg [gof081f - 1 : 0] mt18be0;
reg [DINWIDTH - 1 : 0] tw2f823;
reg [DINWIDTH - 1 : 0] ose08da;
reg [DINWIDTH - 1 : 0] ux23682;
reg [DINWIDTH - 1 : 0] zkda0a2;
reg [DINWIDTH - 1 : 0] aa82893;
reg ba14498;
reg vka24c3;
reg [DINWIDTH - 1 : 0] pu930d4;
reg [DINWIDTH - 1 : 0] czc3511;
reg [DINWIDTH - 1 : 0] uid4469;
reg ria2349;
reg xy11a4a;
reg [DOUTWIDTH - 1 : 0] ho69290;
reg [DOUTWIDTH - 1 : 0] xj4a418;
reg [DOUTWIDTH - 1 : 0] ux9063a;
reg [TAGSWIDTH - 1 : 0] mt18eab;
reg hbc755c;
reg je3aae7;
reg [DOUTWIDTH - 1 : 0] qvab9d3;
reg [DOUTWIDTH - 1 : 0] ipe74e8;
reg [DOUTWIDTH - 1 : 0] gbd3a23;
reg [DOUTWIDTH - 1 : 0] ene88e9;
reg [DOUTWIDTH - 1 : 0] sj23a64;
reg [DOUTWIDTH - 1 : 0] vve992d;
reg [TAGSWIDTH - 1 : 0] hb64b71;
reg [2047:0] vk25b8e;
wire [34:0] fp2dc72;
localparam ld6e396 = 35,hb71cb6 = 32'hfdffc68b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
function [31:0] rv3e73;
input [31:0] value;
for (rv3e73=0; value>0; rv3e73=rv3e73+1) value = value>>1;
endfunction
generate begin : ofc60da   if (INREG == "Enable") begin      if (INSERIAL == "Serial") begin         xy1b553_colorspace #(.psdaa9a     (DINWIDTH      ))         tjaa69b  (.clk            (clk           ),                       .rstn           (rstn          ),                       .ce             (ngb77c            ),                       .sr             (kd5bbe3            ),                       .ph27078            (jc7c771          ),                       .wwc1e36           (pua7f60        ));         su78d89_colorspace #(.psdaa9a     (DINWIDTH      ))         yzb1265      (.clk            (clk           ),                       .rstn           (rstn          ),                       .ce             (ngb77c            ),                       .sr             (kd5bbe3            ),                       .ww4ca1b           (ba14498     ),                       .ph27078            (tw2f823        ),                       .dout0          (gb606af         ),                       .dout1          (aa1abef         ),                       .dout2          (rvafbca         ));      end else begin         xy1b553_colorspace #(.psdaa9a     (DINWIDTH      ))         tjaa69b  (.clk            (clk           ),                       .rstn           (rstn          ),                       .ce             (ngb77c            ),                       .sr             (kd5bbe3            ),                       .ph27078            (jc7c771          ),                       .wwc1e36           (gb606af         ));         xy1b553_colorspace #(.psdaa9a     (DINWIDTH      ))         ho4809c  (.clk            (clk           ),                       .rstn           (rstn          ),                       .ce             (ngb77c            ),                       .sr             (kd5bbe3            ),                       .ph27078            (oh1dc57          ),                       .wwc1e36           (aa1abef         ));         xy1b553_colorspace #(.psdaa9a     (DINWIDTH      ))         yzb18b1  (.clk            (clk           ),                       .rstn           (rstn          ),                       .ce             (ngb77c            ),                       .sr             (kd5bbe3            ),                       .ph27078            (jp715e2          ),                       .wwc1e36           (rvafbca         ));      end   end else begin      if (INSERIAL == "Serial") begin         su78d89_colorspace #(.psdaa9a     (DINWIDTH      ))         yzb1265      (.clk            (clk           ),                       .rstn           (rstn          ),                       .ce             (ngb77c            ),                       .sr             (kd5bbe3            ),                       .ww4ca1b           (ba14498     ),                       .ph27078            (jc7c771          ),                       .dout0          (gb606af         ),                       .dout1          (aa1abef         ),                       .dout2          (rvafbca         ));      end else begin         assign gb606af   = jc7c771;         assign aa1abef   = oh1dc57;         assign rvafbca   = jp715e2;      end   end
end
endgenerate             bnb0774_colorspace #(.TAGSWIDTH       (TAGSWIDTH      ),                     .INSERIAL        (INSERIAL       ),                     .INREG           (INREG          ),                     .LATENCY         (LATENCY-KEEPBLANK))             mrf8dc8 (.tags_in         (jc578b4        ),                     .clk             (clk            ),                     .rstn            (rstn           ),                     .ce              (ngb77c             ),                     .sr              (kd5bbe3             ),                     .inpvalid        (vvddf1d       ),                     .meef2b9       (meef2b9      ),                     .tags_out        (zz1c615     ),                     .ea7de57       (ea7de57      ),                     .outvalid        (gd12433     ));       qg62f86_colorspace # (.CORETYPE         (CORETYPE       ),                    .psdaa9a       (DINWIDTH       ),                    .CWIDTH           (CWIDTH         ),                    .CPOINTS          (CPOINTS        ),                    .ym3b97e     (ym3b97e   ),                    .vk2fc20   (vk2fc20 ),                    .gof081f   (gof081f ),                    .DINSIGN          (DINSIGN        ),                    .INSERIAL         (INSERIAL       ),                    .DEVICE           (DEVICE         ),                    .OPTIMIZE         (OPTIMIZE       ),                    .DSPBLKMULT       (DSPBLKMULT     ),                    .CV_MH            (CV_MH          ),                    .CV_MI            (CV_MI          ),                    .CV_MJ            (CV_MJ          ),                    .CV_MK            (CV_MK          ),                    .CV_NH            (CV_NH          ),                    .CV_NI            (CV_NI          ),                    .CV_NJ            (CV_NJ          ),                    .CV_NK            (CV_NK          ),                    .CV_PH            (CV_PH          ),                    .CV_PI            (CV_PI          ),                    .CV_PJ            (CV_PJ          ),                    .CV_PK            (CV_PK          ))       co24a59 (                    .clk              (clk            ),                    .rstn             (rstn           ),                    .ce               (ngb77c             ),                    .sr               (kd5bbe3             ),                    .meef2b9        (vka24c3      ),                    .din0             (ux23682          ),                    .din1             (zkda0a2          ),                    .din2             (aa82893          ),                    .dout0            (cz51c7a         ),                    .dout1            (th71ea7         ),                    .dout2            (kd7a9fd         ));
         ria7226_colorspace #(                   .yz39132           (gof081f  ),                   .al44ca7    (MSBMETHOD       ),                   .ph329ec    (LSBMETHOD       ),                   .pua7b36         ("Signed"        ),                   .nt3d9b3        (DOUTSIGN        ),                   .ps66cfe        (0               ),                   .CPOINTS          (CPOINTS         ),                   .DOUTPOINTS       (DOUTPOINTS      ),                   .DOUTWIDTH        (DOUTWIDTH       ),                   .ene8af1         (0               ))         dz4578c  (                  .clk               (clk             ),                  .rstn              (rstn            ),                  .ce                (ngb77c              ),                  .sr                (kd5bbe3              ),                  .ph27078               (ale2d18          ),                  .wwc1e36              (hq86704         ));
generate begin : by5248d   if (INSERIAL == "Parallel") begin       ria7226_colorspace #(                  .yz39132            (gof081f  ),                  .al44ca7     (MSBMETHOD       ),                  .ph329ec     (LSBMETHOD       ),                  .pua7b36          ("Signed"        ),                  .nt3d9b3         (DOUTSIGN        ),                  .ps66cfe         (0               ),                  .CPOINTS           (CPOINTS         ),                  .DOUTPOINTS        (DOUTPOINTS      ),                  .DOUTWIDTH         (DOUTWIDTH       ),                  .ene8af1          (0               ))       sj3306d    (                  .clk               (clk             ),                  .rstn              (rstn            ),                  .ce                (ngb77c              ),                  .sr                (kd5bbe3              ),                  .ph27078               (qvb462f          ),                  .wwc1e36              (ba9c11c         ));       ria7226_colorspace #(                  .yz39132            (gof081f  ),                  .al44ca7     (MSBMETHOD       ),                  .ph329ec     (LSBMETHOD       ),                  .pua7b36          ("Signed"        ),                  .nt3d9b3         (DOUTSIGN        ),                  .ps66cfe         (0               ),                  .CPOINTS           (CPOINTS         ),                  .DOUTPOINTS        (DOUTPOINTS      ),                  .DOUTWIDTH         (DOUTWIDTH       ),                  .ene8af1          (0               ))       kq7ded4    (                  .clk               (clk             ),                  .rstn              (rstn            ),                  .ce                (ngb77c              ),                  .sr                (kd5bbe3              ),                  .ph27078               (mt18be0          ),                  .wwc1e36              (ba4718         ));   end
end
if(KEEPBLANK==0) begin   assign outvalid = ria2349;   assign dout0    = ho69290;   assign dout1    = xj4a418;   assign dout2    = ux9063a;   assign tags_out = mt18eab;
end else begin   assign outvalid = hbc755c;   assign dout0    = ene88e9;   assign dout1    = sj23a64;   assign dout2    = vve992d;   assign tags_out = hb64b71;   assign ec9219c = (IOVALID==0) ? 1'b1 : (INSERIAL == "Serial") ? (ria2349 || hbc755c || je3aae7) : (ria2349);   if(DOUTWIDTH>DINWIDTH) begin      assign uk15fae = {pu930d4,{(DOUTWIDTH-DINWIDTH){1'b0}}};      assign rt7eb87 = {czc3511,{(DOUTWIDTH-DINWIDTH){1'b0}}};      assign qvae1f1 = {uid4469,{(DOUTWIDTH-DINWIDTH){1'b0}}};   end else begin      assign uk15fae = pu930d4[DINWIDTH-1:DINWIDTH-DOUTWIDTH];      assign rt7eb87 = czc3511[DINWIDTH-1:DINWIDTH-DOUTWIDTH];      assign qvae1f1 = uid4469[DINWIDTH-1:DINWIDTH-DOUTWIDTH];   end   always @(posedge clk or negedge rstn) begin      if (!rstn) begin         lde30af <= 1'b0;         cb1857e<= 1'b0;         gq87c65    <= {DOUTWIDTH{1'b0}};         byf1941    <= {DOUTWIDTH{1'b0}};         uv6505b    <= {DOUTWIDTH{1'b0}};         ip416ef <= {DOUTWIDTH{1'b0}};      end else if (ngb77c) begin         if (kd5bbe3) begin            lde30af <= 1'b0;            cb1857e<= 1'b0;            gq87c65    <= {DOUTWIDTH{1'b0}};            byf1941    <= {DOUTWIDTH{1'b0}};            uv6505b    <= {DOUTWIDTH{1'b0}};            ip416ef <= {DOUTWIDTH{1'b0}};         end else begin            lde30af <= ria2349;            cb1857e<= hbc755c;            ip416ef <= mt18eab;            if(xy11a4a) begin               gq87c65    <= ho69290;               byf1941    <= xj4a418;               uv6505b    <= ux9063a;            end else begin               gq87c65    <= qvab9d3;               byf1941    <= ipe74e8;               uv6505b    <= gbd3a23;            end         end      end   end      pmi_distributed_shift_reg  #( .pmi_data_width      (3*DINWIDTH ),                                 .pmi_regmode         ("reg"      ),                                 .pmi_shiftreg_type   ("fixed"    ),                                 .pmi_num_shift       (LATENCY-1 ),                                 .pmi_num_width       (je207ce    ),                                                                  .pmi_max_shift       (LATENCY-1 ),                                 .pmi_max_width       (je207ce    ),                                                                  .pmi_init_file       ("none"     ),                                 .pmi_init_file_format("binary"   ),                                 .pmi_family          (DEVICE     ),                                 .module_type         ("pmi_distributed_shift_reg"))   ri2fd71            ( .Din      ({din0,din1,din2}      ),                                 .Addr     ({je207ce{1'b0}}       ),                                 .Clock    (clk                   ),                                 .ClockEn  (ce                    ),                                 .Reset    (~rstn || sr           ),                                 .Q        ({dmcae42,gqb9092,ne42486}));
end
endgenerate
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];vvddf1d<=fp2dc72[2];jc7c771<={din0>>1,fp2dc72[3]};oh1dc57<={din1>>1,fp2dc72[4]};jp715e2<={din2>>1,fp2dc72[5]};jc578b4<={tags_in>>1,fp2dc72[6]};ale2d18<={cz51c7a>>1,fp2dc72[7]};qvb462f<={th71ea7>>1,fp2dc72[8]};mt18be0<={kd7a9fd>>1,fp2dc72[9]};tw2f823<={pua7f60>>1,fp2dc72[10]};ose08da<={offd81a>>1,fp2dc72[11]};ux23682<={gb606af>>1,fp2dc72[12]};zkda0a2<={aa1abef>>1,fp2dc72[13]};aa82893<={rvafbca>>1,fp2dc72[14]};ba14498<=fp2dc72[15];vka24c3<=fp2dc72[16];pu930d4<={dmcae42>>1,fp2dc72[17]};czc3511<={gqb9092>>1,fp2dc72[18]};uid4469<={ne42486>>1,fp2dc72[19]};ria2349<=fp2dc72[20];xy11a4a<=fp2dc72[21];ho69290<={hq86704>>1,fp2dc72[22]};xj4a418<={ba9c11c>>1,fp2dc72[23]};ux9063a<={ba4718>>1,fp2dc72[24]};mt18eab<={zz1c615>>1,fp2dc72[25]};hbc755c<=fp2dc72[26];je3aae7<=fp2dc72[27];qvab9d3<={uk15fae>>1,fp2dc72[28]};ipe74e8<={rt7eb87>>1,fp2dc72[29]};gbd3a23<={qvae1f1>>1,fp2dc72[30]};ene88e9<={gq87c65>>1,fp2dc72[31]};sj23a64<={byf1941>>1,fp2dc72[32]};vve992d<={uv6505b>>1,fp2dc72[33]};hb64b71<={ip416ef>>1,fp2dc72[34]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=inpvalid;vk25b8e[2044]<=din0[0];vk25b8e[2040]<=din1[0];vk25b8e[2032]<=din2[0];vk25b8e[2017]<=tags_in[0];vk25b8e[1987]<=cz51c7a[0];vk25b8e[1963]<=uv6505b[0];vk25b8e[1926]<=th71ea7[0];vk25b8e[1921]<=ba9c11c[0];vk25b8e[1879]<=ip416ef[0];vk25b8e[1805]<=kd7a9fd[0];vk25b8e[1795]<=ba4718[0];vk25b8e[1679]<=meef2b9;vk25b8e[1562]<=pua7f60[0];vk25b8e[1543]<=zz1c615[0];vk25b8e[1310]<=dmcae42[0];vk25b8e[1144]<=ne42486[0];vk25b8e[1076]<=offd81a[0];vk25b8e[1039]<=lde30af;vk25b8e[1023]<=ce;vk25b8e[981]<=byf1941[0];vk25b8e[960]<=hq86704[0];vk25b8e[839]<=ea7de57;vk25b8e[572]<=gqb9092[0];vk25b8e[490]<=gq87c65[0];vk25b8e[480]<=ec9219c;vk25b8e[419]<=rvafbca[0];vk25b8e[245]<=qvae1f1[0];vk25b8e[240]<=gd12433;vk25b8e[209]<=aa1abef[0];vk25b8e[122]<=rt7eb87[0];vk25b8e[104]<=gb606af[0];vk25b8e[61]<=uk15fae[0];vk25b8e[30]<=cb1857e;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module ria7226_colorspace (
              
              clk,
              rstn,
              ce,
              sr,
              ph27078,
              
              wwc1e36
              );
parameter yz39132           = 12;
parameter al44ca7    = "Truncation";
parameter ph329ec    = "Truncation";
parameter pua7b36         = "Unsigned";
parameter nt3d9b3        = "Unsigned";
parameter ps66cfe        = 0;
parameter CPOINTS          = 0;
parameter DOUTPOINTS       = 0;
parameter DOUTWIDTH        = 32;
parameter ene8af1         = 0;
localparam sw212c2 = ((yz39132==DOUTWIDTH && DOUTPOINTS==(ps66cfe+CPOINTS)) && !(pua7b36=="Signed" && nt3d9b3=="Unsigned")) ? 0 : 1;
localparam uxabeb4 = (DOUTPOINTS < ps66cfe+CPOINTS) ? ps66cfe+CPOINTS-DOUTPOINTS : 0;
localparam yx70b70  = 24;
localparam oh85b85 = (pua7b36 == "Unsigned") ? yz39132-uxabeb4 : yz39132-uxabeb4+1;
localparam dz6ed6e = (oh85b85+yx70b70-1)/yx70b70;
localparam fn6eeba = (uxabeb4 == 0 || ph329ec == "Truncation") ? 1 : 0;
localparam hbd75ce = ((al44ca7 == "Truncation") && !(pua7b36 == "Signed" && nt3d9b3 == "Unsigned")) ? 1 : 0;
localparam kqcedb1 = (sw212c2==0) ? 0 :                    (fn6eeba==1 && hbd75ce==1) ? 0 :                    (fn6eeba==1 && hbd75ce==0) ? 1 :                    (fn6eeba==0 && hbd75ce==1) ? dz6ed6e+1 : dz6ed6e+2;
localparam sh6067e = (ene8af1 == 0) ? kqcedb1 : kqcedb1+1;
input                       clk;
input                       rstn;
input                       ce;
input                       sr;
input[yz39132-1:0]           ph27078;
output[DOUTWIDTH-1:0]       wwc1e36;
reg ngb77c;
reg kd5bbe3;
reg [yz39132 - 1 : 0] wy15935;
reg [2047:0] vk25b8e;
wire [2:0] fp2dc72;
localparam ld6e396 = 3,hb71cb6 = 32'hfdffc68b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
 twa8e69_colorspace #(.yz39132         (yz39132       ),        .DOUTWIDTH      (DOUTWIDTH    ),        .sw212c2  (sw212c2),        .ph329ec  (ph329ec),        .al44ca7  (al44ca7),        .yx70b70          (yx70b70        ),        .ps66cfe      (ps66cfe    ),        .CPOINTS        (CPOINTS      ),        .DOUTPOINTS     (DOUTPOINTS   ),        .pua7b36       (pua7b36     ),        .nt3d9b3      (nt3d9b3    ),        .ene8af1       (ene8af1     ))
yz2e0e(        .rstn           (rstn         ),        .clk            (clk          ),        .ce             (ngb77c           ),        .sr             (kd5bbe3           ),        .ph27078            (wy15935          ),        .wwc1e36           (wwc1e36         ));
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];wy15935<={ph27078>>1,fp2dc72[2]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=ph27078[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module bnb0774_colorspace (
               
               clk,                 
               rstn,                
               ce,                  
               sr,                  
               inpvalid,            
               tags_in,             
               tags_out,         
               meef2b9,           
               ea7de57,           
               outvalid             
               );
parameter   TAGSWIDTH        =   8;
parameter   INSERIAL         =   "Serial";
parameter   INREG            =   "Enable";
parameter   LATENCY          =   1;
localparam  dmf474a           =   (INREG == "Enable")? 1 : 0;
input                      clk;
input                      rstn;
input                      ce;
input                      sr;
input                      inpvalid;
input [TAGSWIDTH-1:0]      tags_in;
output                     meef2b9;
output                     ea7de57;
output                     outvalid;
output  [TAGSWIDTH-1:0]    tags_out;
reg  [LATENCY-1:0]         ww68949;
reg  [TAGSWIDTH-1:0]       do25245 [0:LATENCY-1];
integer cm4915d;
reg ngb77c;
reg kd5bbe3;
reg vvddf1d;
reg [TAGSWIDTH - 1 : 0] jc578b4;
reg [LATENCY - 1 : 0] do1e2e8;
reg [2047:0] vk25b8e;
wire [4:0] fp2dc72;
localparam ld6e396 = 5,hb71cb6 = 32'hfdffca8b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
assign outvalid = do1e2e8[LATENCY-1];
generate   if (INSERIAL == "Serial") begin      assign ea7de57 = do1e2e8[1+dmf474a];      assign meef2b9 = do1e2e8[0+dmf474a];   end
endgenerate
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      ww68949   <= {LATENCY{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         ww68949  <= {LATENCY{1'b0}};      end else begin         ww68949  <= {do1e2e8[LATENCY-2:0],vvddf1d};      end   end
end
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      for (cm4915d=0;cm4915d<LATENCY;cm4915d=cm4915d+1) begin         do25245[cm4915d]    <= {{TAGSWIDTH}{1'b0}};      end   end   else if (ngb77c) begin      if (kd5bbe3)  begin         for (cm4915d=0;cm4915d<LATENCY;cm4915d=cm4915d+1) begin            do25245[cm4915d]    <= {{TAGSWIDTH}{1'b0}};         end      end      else begin         do25245[0] <= jc578b4;         for (cm4915d=1;cm4915d<LATENCY;cm4915d=cm4915d+1) begin            do25245[cm4915d]    <= do25245[cm4915d-1];         end      end   end
end
assign tags_out = do25245[LATENCY-1];
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];vvddf1d<=fp2dc72[2];jc578b4<={tags_in>>1,fp2dc72[3]};do1e2e8<={ww68949>>1,fp2dc72[4]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=inpvalid;vk25b8e[2044]<=tags_in[0];vk25b8e[2040]<=ww68949[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module qg62f86_colorspace (
               clk,                 
               rstn,                
               ce,                  
               sr,                  
               meef2b9,           
               din0,                
               din1,                
               din2,                
               dout0,               
               dout1,               
               dout2                
               );
parameter      CORETYPE          = 0;
parameter      psdaa9a        = 12;
parameter      CWIDTH            = 8;
parameter      CPOINTS           =  0;
parameter      ym3b97e      = 20;
parameter      vk2fc20    = 21;
parameter      gof081f    = 22;
parameter      DINSIGN           = "Signed";
parameter      INSERIAL          = "Serial";
parameter      DEVICE            = "ECP2";
parameter      OPTIMIZE          = 0;
parameter      DSPBLKMULT        = "Enable";
parameter      CV_MH             = 0;
parameter      CV_MI             = 0;
parameter      CV_MJ             = 0;
parameter      CV_MK             = 0;
parameter      CV_NH             = 0;
parameter      CV_NI             = 0;
parameter      CV_NJ             = 0;
parameter      CV_NK             = 0;
parameter      CV_PH             = 0;
parameter      CV_PI             = 0;
parameter      CV_PJ             = 0;
parameter      CV_PK             = 0;
input                            clk;
input                            rstn;
input                            ce;
input                            sr;
input                            meef2b9;
input  [psdaa9a-1:0]          din0;
input  [psdaa9a-1:0]          din1;
input  [psdaa9a-1:0]          din2;
output [gof081f-1:0]      dout0;
output [gof081f-1:0]      dout1;
output [gof081f-1:0]      dout2;
reg ngb77c;
reg kd5bbe3;
reg vka24c3;
reg [psdaa9a - 1 : 0] jc7c771;
reg [psdaa9a - 1 : 0] oh1dc57;
reg [psdaa9a - 1 : 0] jp715e2;
reg [2047:0] vk25b8e;
wire [5:0] fp2dc72;
localparam ld6e396 = 6,hb71cb6 = 32'hfdffe06b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
generate begin   if (INSERIAL == "Parallel") begin      if (OPTIMIZE == 0) begin         zm89239_colorspace #(.CORETYPE         (  CORETYPE       ),                           .psdaa9a       (  psdaa9a     ),                           .CWIDTH           (  CWIDTH         ),                           .CPOINTS          (  CPOINTS        ),                           .ym3b97e     (  ym3b97e   ),                           .vk2fc20   (  vk2fc20 ),                           .gof081f   (  gof081f ),                           .DINSIGN          (  DINSIGN        ),                           .DSPBLKMULT       (  DSPBLKMULT     ),                           .INSERIAL         (  INSERIAL   ),                           .DEVICE           (  DEVICE         ),                           .CV_MH            (  CV_MH          ),                           .CV_MI            (  CV_MI          ),                           .CV_MJ            (  CV_MJ          ),                           .CV_MK            (  CV_MK          ),                           .CV_NH            (  CV_NH          ),                           .CV_NI            (  CV_NI          ),                           .CV_NJ            (  CV_NJ          ),                           .CV_NK            (  CV_NK          ),                           .CV_PH            (  CV_PH          ),                           .CV_PI            (  CV_PI          ),                           .CV_PJ            (  CV_PJ          ),                           .CV_PK            (  CV_PK          )                          )         sh41816  (.clk              (  clk            ),                           .rstn             (  rstn           ),                           .ce               (  ngb77c             ),                           .sr               (  kd5bbe3             ),                           .din0             (  jc7c771           ),                           .din1             (  oh1dc57           ),                           .din2             (  jp715e2           ),                           .dout0            (  dout0          ),                           .dout1            (  dout1          ),                           .dout2            (  dout2          )                          );      end else begin         rv6684_colorspace #(.CORETYPE         (  CORETYPE       ),                           .psdaa9a       (  psdaa9a     ),                           .CWIDTH           (  CWIDTH         ),                           .CPOINTS          (  CPOINTS        ),                           .ym3b97e     (  ym3b97e   ),                           .vk2fc20   (  vk2fc20 ),                           .gof081f   (  gof081f ),                           .DINSIGN          (  DINSIGN        ),                           .DSPBLKMULT       (  DSPBLKMULT     ),                           .INSERIAL         (  INSERIAL       ),                           .DEVICE           (  DEVICE         ),                           .CV_MH            (  CV_MH          ),                           .CV_MI            (  CV_MI          ),                           .CV_MJ            (  CV_MJ          ),                           .CV_MK            (  CV_MK          ),                           .CV_NH            (  CV_NH          ),                           .CV_NI            (  CV_NI          ),                           .CV_NJ            (  CV_NJ          ),                           .CV_NK            (  CV_NK          ),                           .CV_PH            (  CV_PH          ),                           .CV_PI            (  CV_PI          ),                           .CV_PJ            (  CV_PJ          ),                           .CV_PK            (  CV_PK          )                          )         sh41816  (.clk              (  clk            ),                           .rstn             (  rstn           ),                           .ce               (  ngb77c             ),                           .sr               (  kd5bbe3             ),                           .din0             (  jc7c771           ),                           .din1             (  oh1dc57           ),                           .din2             (  jp715e2           ),                           .dout0            (  dout0          ),                           .dout1            (  dout1          ),                           .dout2            (  dout2          )                          );      end   end else begin      pf6b769_colorspace #(.CORETYPE         (  CORETYPE       ),                        .psdaa9a       (  psdaa9a     ),                        .CWIDTH           (  CWIDTH         ),                        .CPOINTS          (  CPOINTS        ),                        .ym3b97e     (  ym3b97e   ),                        .vk2fc20   (  vk2fc20 ),                        .gof081f   (  gof081f ),                        .DINSIGN          (  DINSIGN        ),                        .DSPBLKMULT       (  DSPBLKMULT     ),                        .INSERIAL         (  INSERIAL       ),                        .DEVICE           (  DEVICE         ),                        .CV_MH            (  CV_MH          ),                        .CV_MI            (  CV_MI          ),                        .CV_MJ            (  CV_MJ          ),                        .CV_MK            (  CV_MK          ),                        .CV_NH            (  CV_NH          ),                        .CV_NI            (  CV_NI          ),                        .CV_NJ            (  CV_NJ          ),                        .CV_NK            (  CV_NK          ),                        .CV_PH            (  CV_PH          ),                        .CV_PI            (  CV_PI          ),                        .CV_PJ            (  CV_PJ          ),                        .CV_PK            (  CV_PK          )                       )      hoe4c89  (.clk              (  clk            ),                        .rstn             (  rstn           ),                        .ce               (  ngb77c             ),                        .sr               (  kd5bbe3             ),                        .meef2b9        (  vka24c3      ),                        .din0             (  jc7c771           ),                        .din1             (  oh1dc57           ),                        .din2             (  jp715e2           ),                        .dout0            (  dout0          )                       );   end
end
endgenerate
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];vka24c3<=fp2dc72[2];jc7c771<={din0>>1,fp2dc72[3]};oh1dc57<={din1>>1,fp2dc72[4]};jp715e2<={din2>>1,fp2dc72[5]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=meef2b9;vk25b8e[2044]<=din0[0];vk25b8e[2041]<=din1[0];vk25b8e[2034]<=din2[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module gbe8249_colorspace (
               rstn,
               clk,
               ce,
               sr,
               jc4d981,
               dm6cc0b,
               wwc1e36
            );
parameter   yz39132   = 32;
parameter   bn81692    = "Unsigned";
parameter   yx70b70    = 16;
localparam  fn5a4b3     = 1'b1;
localparam  dzd259e    = 1'b0;
localparam  gq92cf6   = yz39132+1;
localparam  cob3d8a     = (yz39132+yx70b70-1)/yx70b70;
localparam  ux8a1fc    = yz39132%yx70b70;
input                   rstn;
input                   clk;
input                   ce;
input                   sr;
input [yz39132-1:0]      jc4d981;
input [yz39132-1:0]      dm6cc0b;
output[gq92cf6-1:0]      wwc1e36;
wire[yx70b70*cob3d8a-1:0]    db22692;
wire[yx70b70*cob3d8a-1:0]    nrd25b4;
genvar ie92da6,zm96d31,ecb698b;
reg             gdb4c58[0:cob3d8a] ;
wire[yx70b70-1:0] bn8b140[0:cob3d8a-1];
wire[yx70b70-1:0] zz281d2[0:cob3d8a-1];
reg [yx70b70-1:0] vk3a5fd[0:cob3d8a-1][0:cob3d8a-1] ;
reg [yx70b70-1:0] wjfd7ce[0:cob3d8a-1][0:cob3d8a-1] ;
reg [yx70b70-1:0] goce8f7[0:cob3d8a-1][0:cob3d8a-1] ;
reg ngb77c;
reg kd5bbe3;
reg [yz39132 - 1 : 0] yxc62eb;
reg [yz39132 - 1 : 0] jr8bae8;
reg [yx70b70 * cob3d8a - 1 : 0] tu5d19b;
reg [yx70b70 * cob3d8a - 1 : 0] wl336e1;
reg [2047:0] vk25b8e;
wire [5:0] fp2dc72;
localparam ld6e396 = 6,hb71cb6 = 32'hfdffca8b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
assign db22692 = ux8a1fc==0 ? yxc62eb : bn81692=="Signed" ? {{(yx70b70-ux8a1fc){yxc62eb[yz39132-1]}},yxc62eb}:                                {{(yx70b70-ux8a1fc){dzd259e}},yxc62eb};
assign nrd25b4 = ux8a1fc==0 ? jr8bae8 : bn81692=="Signed" ? {{(yx70b70-ux8a1fc){jr8bae8[yz39132-1]}},jr8bae8}:                                {{(yx70b70-ux8a1fc){dzd259e}},jr8bae8};
generate
begin   for (ie92da6=0;ie92da6<cob3d8a;ie92da6=ie92da6+1) begin:rg57f29      assign bn8b140[ie92da6] = tu5d19b[yx70b70*(ie92da6+1)-1:yx70b70*ie92da6];      assign zz281d2[ie92da6] = wl336e1[yx70b70*(ie92da6+1)-1:yx70b70*ie92da6];      for (zm96d31=0;zm96d31<ie92da6;zm96d31=zm96d31+1) begin:mgbc097         always @(posedge clk or negedge rstn)         begin            if (rstn == dzd259e) begin               vk3a5fd[ie92da6][zm96d31] <= {yx70b70{dzd259e}};               wjfd7ce[ie92da6][zm96d31] <= {yx70b70{dzd259e}};            end else if (ngb77c == fn5a4b3) begin               if (kd5bbe3) begin                  vk3a5fd[ie92da6][zm96d31] <= {yx70b70{dzd259e}};                  wjfd7ce[ie92da6][zm96d31] <= {yx70b70{dzd259e}};               end else begin                  vk3a5fd[ie92da6][zm96d31] <= zm96d31==0 ? bn8b140[ie92da6] : vk3a5fd[ie92da6][zm96d31-1];                  wjfd7ce[ie92da6][zm96d31] <= zm96d31==0 ? zz281d2[ie92da6] : wjfd7ce[ie92da6][zm96d31-1];               end            end         end      end      if (ie92da6 == cob3d8a-1) begin         always @(posedge clk or negedge rstn)         begin            if (rstn == dzd259e)               {gdb4c58[ie92da6],goce8f7[ie92da6][ie92da6]} <= {(yx70b70+1){dzd259e}};            else if (ngb77c == fn5a4b3) begin               if (kd5bbe3 == fn5a4b3)                  {gdb4c58[ie92da6],goce8f7[ie92da6][ie92da6]} <= {(yx70b70+1){dzd259e}};               else if (bn81692 == "Unsigned")                  {gdb4c58[ie92da6],goce8f7[ie92da6][ie92da6]} <= ie92da6==0 ?  bn8b140[0]+zz281d2[0]+1'b0 :                              vk3a5fd[ie92da6][ie92da6-1]+wjfd7ce[ie92da6][ie92da6-1]+gdb4c58[ie92da6-1];               else                  {gdb4c58[ie92da6],goce8f7[ie92da6][ie92da6]} <= ie92da6==0 ?  {bn8b140[0][yx70b70-1],bn8b140[0]}+{zz281d2[0][yx70b70-1],zz281d2[0]}+1'b0 :                              {vk3a5fd[ie92da6][ie92da6-1][yx70b70-1],vk3a5fd[ie92da6][ie92da6-1]}+{wjfd7ce[ie92da6][ie92da6-1][yx70b70-1],wjfd7ce[ie92da6][ie92da6-1]}+gdb4c58[ie92da6-1];            end         end      end else begin         always @(posedge clk or negedge rstn)         begin            if (rstn == dzd259e)               {gdb4c58[ie92da6],goce8f7[ie92da6][ie92da6]} <= {(yx70b70+1){dzd259e}};            else if (ngb77c == fn5a4b3) begin               if (kd5bbe3 == fn5a4b3)                  {gdb4c58[ie92da6],goce8f7[ie92da6][ie92da6]} <= {(yx70b70+1){dzd259e}};               else                  {gdb4c58[ie92da6],goce8f7[ie92da6][ie92da6]} <= ie92da6==0 ?  bn8b140[0]+zz281d2[0]+1'b0 :                           vk3a5fd[ie92da6][ie92da6-1]+wjfd7ce[ie92da6][ie92da6-1]+gdb4c58[ie92da6-1];            end         end      end      for (zm96d31=ie92da6+1;zm96d31<cob3d8a;zm96d31=zm96d31+1) begin:kf1d7c4         always @(posedge clk or negedge rstn)         begin            if (rstn == dzd259e)               goce8f7[ie92da6][zm96d31] <= {(yx70b70+1){dzd259e}};            else if (ngb77c == fn5a4b3) begin               if (kd5bbe3 == fn5a4b3)                  goce8f7[ie92da6][zm96d31] <= {(yx70b70+1){dzd259e}};               else                  goce8f7[ie92da6][zm96d31] <= goce8f7[ie92da6][zm96d31-1];            end         end      end   end   if (ux8a1fc == 0) begin      for (ie92da6=0;ie92da6<cob3d8a;ie92da6=ie92da6+1) begin:ux2323e         assign wwc1e36[yx70b70*(ie92da6+1)-1:yx70b70*ie92da6] = goce8f7[ie92da6][cob3d8a-1];      end      assign wwc1e36[gq92cf6-1] = gdb4c58[cob3d8a-1];   end else begin      for (ie92da6=0;ie92da6<cob3d8a-1;ie92da6=ie92da6+1) begin:ux85312         assign wwc1e36[yx70b70*(ie92da6+1)-1:yx70b70*ie92da6] = goce8f7[ie92da6][cob3d8a-1];      end      assign wwc1e36[gq92cf6-1:gq92cf6-ux8a1fc-1] = goce8f7[cob3d8a-1][cob3d8a-1][ux8a1fc:0];   end
end
endgenerate
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];yxc62eb<={jc4d981>>1,fp2dc72[2]};jr8bae8<={dm6cc0b>>1,fp2dc72[3]};tu5d19b<={db22692>>1,fp2dc72[4]};wl336e1<={nrd25b4>>1,fp2dc72[5]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=jc4d981[0];vk25b8e[2044]<=dm6cc0b[0];vk25b8e[2040]<=db22692[0];vk25b8e[2032]<=nrd25b4[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module zm89239_colorspace (
                     clk,   
                     rstn,
                     ce,
                     sr,
                     din0,
                     din1,
                     din2,
                     dout0,
                     dout1,
                     dout2);
parameter      CORETYPE          = 0;
parameter      psdaa9a        = 12;
parameter      CWIDTH            = 8;
parameter      CPOINTS           = 0;
parameter      ym3b97e      = 20;
parameter      vk2fc20    = 21;
parameter      gof081f    = 22;
parameter      DINSIGN           = "Signed";
parameter      DSPBLKMULT        = "Enable";
parameter      INSERIAL          = "Serial";
parameter      DEVICE            = "ECP2";
parameter      CV_MH             = 0;
parameter      CV_MI             = 0;
parameter      CV_MJ             = 0;
parameter      CV_MK             = 0;
parameter      CV_NH             = 0;
parameter      CV_NI             = 0;
parameter      CV_NJ             = 0;
parameter      CV_NK             = 0;
parameter      CV_PH             = 0;
parameter      CV_PI             = 0;
parameter      CV_PJ             = 0;
parameter      CV_PK             = 0;
localparam     qiadca             =  DINSIGN == "Signed" ? 1'b1 : 1'b0;
input                         clk;
input                         rstn;
input                         ce;
input                         sr;
input  [psdaa9a-1:0]       din0;
input  [psdaa9a-1:0]       din1;
input  [psdaa9a-1:0]       din2;
output [gof081f-1:0]   dout0;
output [gof081f-1:0]   dout1;
output [gof081f-1:0]   dout2;
wire   [psdaa9a-1:0]       czfd6b8 [0:2];
wire   [CWIDTH-1:0]           th5ae22 [0:2][0:2];
wire   [ym3b97e-1:0]     zmb88be [0:2];
wire   [ym3b97e-1:0]     nt22f98 [0:2][0:2];
wire   [ym3b97e-1:0]     irbe63d [0:2][0:2];
wire   [vk2fc20-1:0]   ou98f6f;
reg    [ym3b97e-1:0]     fp3dbc6 [0:2][0:2];
reg    [vk2fc20-1:0]   qt6f1bc [0:2];
reg    [vk2fc20-1:0]   wjc6f21 [0:2];
reg    [gof081f-1:0]   aabc866 [0:2];
reg    [psdaa9a-1:0]       ym2198b;
reg    [psdaa9a-1:0]       ho662c7;
reg    [psdaa9a-1:0]       fp8b1d0;
genvar zm96d31,ecb698b;
reg ngb77c;
reg kd5bbe3;
reg [psdaa9a - 1 : 0] jc7c771;
reg [psdaa9a - 1 : 0] oh1dc57;
reg [psdaa9a - 1 : 0] jp715e2;
reg [vk2fc20 - 1 : 0] ui56a8c;
reg [psdaa9a - 1 : 0] xlaa30e;
reg [psdaa9a - 1 : 0] tw8c3b4;
reg [psdaa9a - 1 : 0] pued16;
reg [2047:0] vk25b8e;
wire [8:0] fp2dc72;
localparam ld6e396 = 9,hb71cb6 = 32'hfdffd42b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
generate begin : ou97931   assign zmb88be[0]    = CV_MK;   assign zmb88be[1]    = CV_NK;   assign zmb88be[2]    = CV_PK;   assign th5ae22[0][0] = CV_MH ;   assign th5ae22[0][1] = CV_MI ;   assign th5ae22[0][2] = CV_MJ ;   assign th5ae22[1][0] = CV_NH ;   assign th5ae22[1][1] = CV_NI ;   assign th5ae22[1][2] = CV_NJ ;   assign th5ae22[2][0] = CV_PH ;   assign th5ae22[2][1] = CV_PI ;   assign th5ae22[2][2] = CV_PJ ;   assign czfd6b8[0]    =  jc7c771;   assign czfd6b8[1]    =  oh1dc57;   assign czfd6b8[2]    =  jp715e2;   for (zm96d31=0;zm96d31<3;zm96d31=zm96d31+1) begin : gq2e522      for (ecb698b=0;ecb698b<3;ecb698b=ecb698b+1) begin : qi101ae            if (DSPBLKMULT == "Enable") begin             pmi_dsp_mult   #(.pmi_dataa_width           (psdaa9a    ),                              .pmi_datab_width           (CWIDTH         ),                              .pmi_additional_pipeline   (1              ),                              .pmi_input_reg             ("on"           ),                              .pmi_output_reg            ("on"           ),                              .pmi_family                (DEVICE         ),                              .pmi_gsr                   ("enable"       ),                              .pmi_source_control_a      ("parallel"     ),                              .pmi_source_control_b      ("parallel"     ),                              .pmi_reg_inputa_clk        ("CLK0"         ),                              .pmi_reg_inputa_ce         ("CE0"          ),                              .pmi_reg_inputa_rst        ("RST0"         ),                              .pmi_reg_inputb_clk        ("CLK0"         ),                              .pmi_reg_inputb_ce         ("CE0"          ),                              .pmi_reg_inputb_rst        ("RST0"         ),                              .pmi_reg_pipeline_clk      ("CLK0"         ),                              .pmi_reg_pipeline_ce       ("CE0"          ),                              .pmi_reg_pipeline_rst      ("RST0"         ),                              .pmi_reg_output_clk        ("CLK0"         ),                              .pmi_reg_output_ce         ("CE0"          ),                              .pmi_reg_output_rst        ("RST0"         ),                              .pmi_reg_signeda_clk       ("CLK0"         ),                              .pmi_reg_signeda_ce        ("CE0"          ),                              .pmi_reg_signeda_rst       ("RST0"         ),                              .pmi_reg_signedb_clk       ("CLK0"         ),                              .pmi_reg_signedb_ce        ("CE0"          ),                              .pmi_reg_signedb_rst       ("RST0"         ),                              .pmi_pipelined_mode        ("off"          ),                              .module_type               ("pmi_dsp_mult" )                              )              xj71b9c (                              .A                         (czfd6b8[ecb698b]         ),                              .B                         (th5ae22[zm96d31][ecb698b]     ),                              .SRIA                      (               ),                              .SRIB                      (               ),                              .CLK0                      (clk            ),                              .CLK1                      (clk            ),                              .CLK2                      (clk            ),                              .CLK3                      (clk            ),                              .CE0                       (ce             ),                              .CE1                       (ce             ),                              .CE2                       (ce             ),                              .CE3                       (ce             ),                              .RST0                      (~rstn          ),                              .RST1                      (~rstn          ),                              .RST2                      (~rstn          ),                              .RST3                      (~rstn          ),                              .SignA                     (qiadca          ),                              .SignB                     (1'b1           ),                              .SourceA                   (1'b0           ),                              .SourceB                   (1'b0           ),                              .P                         (nt22f98[zm96d31][ecb698b]),                              .SROA                      (               ),                              .SROB                      (               ));               assign irbe63d[zm96d31][ecb698b] = nt22f98[zm96d31][ecb698b][ym3b97e-1:0];            end else begin                  always @(posedge clk or negedge rstn) begin                      if (!rstn) begin                         fp3dbc6[zm96d31][ecb698b] <= {ym3b97e{1'b0}};                      end else if (ngb77c) begin                         if (kd5bbe3) begin                            fp3dbc6[zm96d31][ecb698b] <= {ym3b97e{1'b0}};                         end else begin                            fp3dbc6[zm96d31][ecb698b] <= nt22f98[zm96d31][ecb698b];                         end                      end                   end                     db199ce_colorspace # (.psdaa9a                (psdaa9a          ),                              .sj39da8                 (CWIDTH              ),                              .jc76a28                     (DINSIGN             ),                              .lsa8a16                     ("Signed"            ))                    hb450b2  (.clk                       (clk                 ),                              .rstn                      (rstn                ),                              .ce                        (ngb77c                  ),                              .sr                        (kd5bbe3                  ),                              .pub26f4                  (czfd6b8[ecb698b]              ),                              .uide8d7                  (th5ae22[zm96d31][ecb698b]          ),                              .irbe63d                  (nt22f98[zm96d31][ecb698b]   ));                    assign irbe63d[zm96d31][ecb698b] = fp3dbc6[zm96d31][ecb698b][ym3b97e-1:0];            end      end   end
end
endgenerate
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      ym2198b <= {psdaa9a{1'b0}};      ho662c7 <= {psdaa9a{1'b0}};      fp8b1d0  <= {psdaa9a{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         ym2198b <= {psdaa9a{1'b0}};         ho662c7 <= {psdaa9a{1'b0}};         fp8b1d0  <= {psdaa9a{1'b0}};      end else begin         ym2198b <= jc7c771;         ho662c7 <= xlaa30e;         fp8b1d0  <= tw8c3b4;      end   end
end
generate begin : uv65b53   if (CPOINTS == 0) begin      if (DINSIGN == "Signed") begin        assign ou98f6f   =  {{(vk2fc20-psdaa9a-CPOINTS){pued16[psdaa9a-1]}},pued16};      end else begin        assign ou98f6f   =  {{(vk2fc20-psdaa9a-CPOINTS){1'b0}},pued16};      end   end else begin      if (DINSIGN == "Signed") begin        assign ou98f6f   =  {{(vk2fc20-psdaa9a-CPOINTS){pued16[psdaa9a-1]}},pued16,{CPOINTS{1'b0}}};      end else begin        assign ou98f6f   =  {{(vk2fc20-psdaa9a-CPOINTS){1'b0}},pued16,{CPOINTS{1'b0}}};      end   end   if (CORETYPE == 0 || CORETYPE == 1 || CORETYPE == 2 || CORETYPE == 3 || CORETYPE == 4) begin      always @(posedge clk or negedge rstn) begin         if (!rstn) begin            qt6f1bc[0] <= {vk2fc20{1'b0}} ;            wjc6f21[0] <= {vk2fc20{1'b0}} ;            aabc866[0] <= {gof081f{1'b0}} ;            qt6f1bc[1] <= {vk2fc20{1'b0}} ;            wjc6f21[1] <= {vk2fc20{1'b0}} ;            aabc866[1] <= {gof081f{1'b0}} ;            qt6f1bc[2] <= {vk2fc20{1'b0}} ;            wjc6f21[2] <= {vk2fc20{1'b0}} ;            aabc866[2] <= {gof081f{1'b0}} ;         end else if (ngb77c) begin            if (kd5bbe3) begin               qt6f1bc[0] <= {vk2fc20{1'b0}} ;               wjc6f21[0] <= {vk2fc20{1'b0}} ;               aabc866[0] <= {gof081f{1'b0}} ;               qt6f1bc[1] <= {vk2fc20{1'b0}} ;               wjc6f21[1] <= {vk2fc20{1'b0}} ;               aabc866[1] <= {gof081f{1'b0}} ;               qt6f1bc[2] <= {vk2fc20{1'b0}} ;               wjc6f21[2] <= {vk2fc20{1'b0}} ;               aabc866[2] <= {gof081f{1'b0}} ;            end else begin               qt6f1bc[0] <= {irbe63d[0][0][ym3b97e-1],irbe63d[0][0]} + {irbe63d[0][1][ym3b97e-1],irbe63d[0][1]};               wjc6f21[0] <= {irbe63d[0][2][ym3b97e-1],irbe63d[0][2]} + {zmb88be[0][ym3b97e-1],zmb88be[0]} ;               aabc866[0] <= {qt6f1bc[0][vk2fc20-1],qt6f1bc[0]}     + {wjc6f21[0][vk2fc20-1],wjc6f21[0]};               qt6f1bc[1] <= {irbe63d[1][0][ym3b97e-1],irbe63d[1][0]} + {irbe63d[1][1][ym3b97e-1],irbe63d[1][1]};               wjc6f21[1] <= {irbe63d[1][2][ym3b97e-1],irbe63d[1][2]} + {zmb88be[1][ym3b97e-1],zmb88be[1]} ;               aabc866[1] <= {qt6f1bc[1][vk2fc20-1],qt6f1bc[1]}     + {wjc6f21[1][vk2fc20-1],wjc6f21[1]};               qt6f1bc[2] <= {irbe63d[2][0][ym3b97e-1],irbe63d[2][0]} + {irbe63d[2][1][ym3b97e-1],irbe63d[2][1]};               wjc6f21[2] <= {irbe63d[2][2][ym3b97e-1],irbe63d[2][2]} + {zmb88be[2][ym3b97e-1],zmb88be[2]} ;               aabc866[2] <= {qt6f1bc[2][vk2fc20-1],qt6f1bc[2]}     + {wjc6f21[2][vk2fc20-1],wjc6f21[2]};            end         end      end   end else if (CORETYPE == 5 || CORETYPE == 6) begin      always @(posedge clk or negedge rstn) begin         if (!rstn) begin            qt6f1bc[0] <= {vk2fc20{1'b0}} ;            wjc6f21[0] <= {vk2fc20{1'b0}} ;            aabc866[0] <= {gof081f{1'b0}} ;            qt6f1bc[1] <= {vk2fc20{1'b0}} ;            wjc6f21[1] <= {vk2fc20{1'b0}} ;            aabc866[1] <= {gof081f{1'b0}} ;            qt6f1bc[2] <= {vk2fc20{1'b0}} ;            wjc6f21[2] <= {vk2fc20{1'b0}} ;            aabc866[2] <= {gof081f{1'b0}} ;         end else if (ngb77c) begin            if (kd5bbe3) begin               qt6f1bc[0] <= {vk2fc20{1'b0}} ;               wjc6f21[0] <= {vk2fc20{1'b0}} ;               aabc866[0] <= {gof081f{1'b0}} ;               qt6f1bc[1] <= {vk2fc20{1'b0}} ;               wjc6f21[1] <= {vk2fc20{1'b0}} ;               aabc866[1] <= {gof081f{1'b0}} ;               qt6f1bc[2] <= {vk2fc20{1'b0}} ;               wjc6f21[2] <= {vk2fc20{1'b0}} ;               aabc866[2] <= {gof081f{1'b0}} ;            end else begin               qt6f1bc[0] <= {irbe63d[0][0][ym3b97e-1],irbe63d[0][0]};               wjc6f21[0] <= {irbe63d[0][2][ym3b97e-1],irbe63d[0][2]} + {zmb88be[0][ym3b97e-1],zmb88be[0]} ;               aabc866[0] <= {qt6f1bc[0][vk2fc20-1],qt6f1bc[0]}     + {wjc6f21[0][vk2fc20-1],wjc6f21[0]};               qt6f1bc[1] <= {irbe63d[0][0][ym3b97e-1],irbe63d[0][0]} + {irbe63d[1][1][ym3b97e-1],irbe63d[1][1]};               wjc6f21[1] <= {irbe63d[1][2][ym3b97e-1],irbe63d[1][2]} + {zmb88be[1][ym3b97e-1],zmb88be[1]} ;               aabc866[1] <= {qt6f1bc[1][vk2fc20-1],qt6f1bc[1]}     + {wjc6f21[1][vk2fc20-1],wjc6f21[1]};               qt6f1bc[2] <= {irbe63d[0][0][ym3b97e-1],irbe63d[0][0]} + {irbe63d[2][1][ym3b97e-1],irbe63d[2][1]};               wjc6f21[2] <= {zmb88be[2][ym3b97e-1],zmb88be[2]} ;               aabc866[2] <= {qt6f1bc[2][vk2fc20-1],qt6f1bc[2]}     + {wjc6f21[2][vk2fc20-1],wjc6f21[2]};            end         end      end   end else if (CORETYPE == 7 || CORETYPE == 8) begin      always @(posedge clk or negedge rstn) begin         if (!rstn) begin            qt6f1bc[0] <= {vk2fc20{1'b0}} ;            wjc6f21[0] <= {vk2fc20{1'b0}} ;            aabc866[0] <= {gof081f{1'b0}} ;            qt6f1bc[1] <= {vk2fc20{1'b0}} ;            wjc6f21[1] <= {vk2fc20{1'b0}} ;            aabc866[1] <= {gof081f{1'b0}} ;            qt6f1bc[2] <= {vk2fc20{1'b0}} ;            wjc6f21[2] <= {vk2fc20{1'b0}} ;            aabc866[2] <= {gof081f{1'b0}} ;         end else if (ngb77c) begin            if (kd5bbe3) begin               qt6f1bc[0] <= {vk2fc20{1'b0}} ;               wjc6f21[0] <= {vk2fc20{1'b0}} ;               aabc866[0] <= {gof081f{1'b0}} ;               qt6f1bc[1] <= {vk2fc20{1'b0}} ;               wjc6f21[1] <= {vk2fc20{1'b0}} ;               aabc866[1] <= {gof081f{1'b0}} ;               qt6f1bc[2] <= {vk2fc20{1'b0}} ;               wjc6f21[2] <= {vk2fc20{1'b0}} ;               aabc866[2] <= {gof081f{1'b0}} ;            end else begin               qt6f1bc[0] <= ui56a8c;               wjc6f21[0] <= {irbe63d[0][2][ym3b97e-1],irbe63d[0][2]} + {zmb88be[0][ym3b97e-1],zmb88be[0]} ;               aabc866[0] <= {qt6f1bc[0][vk2fc20-1],qt6f1bc[0]}     + {wjc6f21[0][vk2fc20-1],wjc6f21[0]};
               qt6f1bc[1] <= ui56a8c + {irbe63d[1][1][ym3b97e-1],irbe63d[1][1]};               wjc6f21[1] <= {irbe63d[1][2][ym3b97e-1],irbe63d[1][2]} + {zmb88be[1][ym3b97e-1],zmb88be[1]} ;               aabc866[1] <= {qt6f1bc[1][vk2fc20-1],qt6f1bc[1]}     + {wjc6f21[1][vk2fc20-1],wjc6f21[1]};               qt6f1bc[2] <= ui56a8c + {irbe63d[2][1][ym3b97e-1],irbe63d[2][1]};               wjc6f21[2] <= {zmb88be[2][ym3b97e-1],zmb88be[2]};               aabc866[2] <= {qt6f1bc[2][vk2fc20-1],qt6f1bc[2]}     + {wjc6f21[2][vk2fc20-1],wjc6f21[2]};            end         end      end   end else if (CORETYPE == 9) begin       always @(posedge clk or negedge rstn) begin         if (!rstn) begin            qt6f1bc[0] <= {vk2fc20{1'b0}} ;            wjc6f21[0] <= {vk2fc20{1'b0}} ;            aabc866[0] <= {gof081f{1'b0}} ;            qt6f1bc[1] <= {vk2fc20{1'b0}} ;            wjc6f21[1] <= {vk2fc20{1'b0}} ;            aabc866[1] <= {gof081f{1'b0}} ;            qt6f1bc[2] <= {vk2fc20{1'b0}} ;            wjc6f21[2] <= {vk2fc20{1'b0}} ;            aabc866[2] <= {gof081f{1'b0}} ;         end else if (ngb77c) begin            if (kd5bbe3) begin               qt6f1bc[0] <= {vk2fc20{1'b0}} ;               wjc6f21[0] <= {vk2fc20{1'b0}} ;               aabc866[0] <= {gof081f{1'b0}} ;               qt6f1bc[1] <= {vk2fc20{1'b0}} ;               wjc6f21[1] <= {vk2fc20{1'b0}} ;               aabc866[1] <= {gof081f{1'b0}} ;               qt6f1bc[2] <= {vk2fc20{1'b0}} ;               wjc6f21[2] <= {vk2fc20{1'b0}} ;               aabc866[2] <= {gof081f{1'b0}} ;            end else begin               qt6f1bc[0] <=  ui56a8c;               wjc6f21[0] <=  {irbe63d[0][2][ym3b97e-1],irbe63d[0][2]};               aabc866[0] <=  {qt6f1bc[0][vk2fc20-1],qt6f1bc[0]}     + {wjc6f21[0][vk2fc20-1],wjc6f21[0]};
               qt6f1bc[1] <=  ui56a8c;               wjc6f21[1] <=  {irbe63d[1][1][ym3b97e-1],irbe63d[1][1]} + {irbe63d[1][2][ym3b97e-1],irbe63d[1][2]};               aabc866[1] <=  {qt6f1bc[1][vk2fc20-1],qt6f1bc[1]}     + {wjc6f21[1][vk2fc20-1],wjc6f21[1]};               qt6f1bc[2] <=  ui56a8c;               wjc6f21[2] <=  {irbe63d[2][1][ym3b97e-1],irbe63d[2][1]};               aabc866[2] <=  {qt6f1bc[2][vk2fc20-1],qt6f1bc[2]}     + {wjc6f21[2][vk2fc20-1],wjc6f21[2]};            end         end      end   end else if (CORETYPE == 10 || CORETYPE == 12) begin      always @(posedge clk or negedge rstn) begin         if (!rstn) begin            qt6f1bc[0] <= {vk2fc20{1'b0}} ;            wjc6f21[0] <= {vk2fc20{1'b0}} ;            aabc866[0] <= {gof081f{1'b0}} ;            qt6f1bc[1] <= {vk2fc20{1'b0}} ;            wjc6f21[1] <= {vk2fc20{1'b0}} ;            aabc866[1] <= {gof081f{1'b0}} ;            qt6f1bc[2] <= {vk2fc20{1'b0}} ;            wjc6f21[2] <= {vk2fc20{1'b0}} ;            aabc866[2] <= {gof081f{1'b0}} ;         end else if (ngb77c) begin            if (kd5bbe3) begin               qt6f1bc[0] <= {vk2fc20{1'b0}} ;               wjc6f21[0] <= {vk2fc20{1'b0}} ;               aabc866[0] <= {gof081f{1'b0}} ;               qt6f1bc[1] <= {vk2fc20{1'b0}} ;               wjc6f21[1] <= {vk2fc20{1'b0}} ;               aabc866[1] <= {gof081f{1'b0}} ;               qt6f1bc[2] <= {vk2fc20{1'b0}} ;               wjc6f21[2] <= {vk2fc20{1'b0}} ;               aabc866[2] <= {gof081f{1'b0}} ;            end else begin               qt6f1bc[0] <=  {irbe63d[0][0][ym3b97e-1],irbe63d[0][0]} + {irbe63d[0][1][ym3b97e-1],irbe63d[0][1]};               wjc6f21[0] <=  {irbe63d[0][2][ym3b97e-1],irbe63d[0][2]};               aabc866[0] <=  {qt6f1bc[0][vk2fc20-1],qt6f1bc[0]}     + {wjc6f21[0][vk2fc20-1],wjc6f21[0]};
               qt6f1bc[1] <=  {irbe63d[1][0][ym3b97e-1],irbe63d[1][0]} + {irbe63d[1][1][ym3b97e-1],irbe63d[1][1]};               wjc6f21[1] <=  {irbe63d[1][2][ym3b97e-1],irbe63d[1][2]};               aabc866[1] <=  {qt6f1bc[1][vk2fc20-1],qt6f1bc[1]}     + {wjc6f21[1][vk2fc20-1],wjc6f21[1]};
               qt6f1bc[2] <=  {irbe63d[2][0][ym3b97e-1],irbe63d[2][0]} + {irbe63d[2][1][ym3b97e-1],irbe63d[2][1]};               wjc6f21[2] <=  {irbe63d[2][2][ym3b97e-1],irbe63d[2][2]};               aabc866[2] <=  {qt6f1bc[2][vk2fc20-1],qt6f1bc[2]}     + {wjc6f21[2][vk2fc20-1],wjc6f21[2]};            end         end      end   end else if (CORETYPE == 11) begin       always @(posedge clk or negedge rstn) begin         if (!rstn) begin            qt6f1bc[0] <= {vk2fc20{1'b0}} ;            wjc6f21[0] <= {vk2fc20{1'b0}} ;            aabc866[0] <= {gof081f{1'b0}} ;            qt6f1bc[1] <= {vk2fc20{1'b0}} ;            wjc6f21[1] <= {vk2fc20{1'b0}} ;            aabc866[1] <= {gof081f{1'b0}} ;            qt6f1bc[2] <= {vk2fc20{1'b0}} ;            wjc6f21[2] <= {vk2fc20{1'b0}} ;            aabc866[2] <= {gof081f{1'b0}} ;         end else if (ngb77c) begin            if (kd5bbe3) begin               qt6f1bc[0] <= {vk2fc20{1'b0}} ;               wjc6f21[0] <= {vk2fc20{1'b0}} ;               aabc866[0] <= {gof081f{1'b0}} ;               qt6f1bc[1] <= {vk2fc20{1'b0}} ;               wjc6f21[1] <= {vk2fc20{1'b0}} ;               aabc866[1] <= {gof081f{1'b0}} ;               qt6f1bc[2] <= {vk2fc20{1'b0}} ;               wjc6f21[2] <= {vk2fc20{1'b0}} ;               aabc866[2] <= {gof081f{1'b0}} ;            end else begin               qt6f1bc[0] <=  ui56a8c;               wjc6f21[0] <=  {irbe63d[0][1][ym3b97e-1],irbe63d[0][1]} + {irbe63d[0][2][ym3b97e-1],irbe63d[0][2]};               aabc866[0] <=  {qt6f1bc[0][vk2fc20-1],qt6f1bc[0]}     + {wjc6f21[0][vk2fc20-1],wjc6f21[0]};
               qt6f1bc[1] <=  ui56a8c;               wjc6f21[1] <=  {irbe63d[1][1][ym3b97e-1],irbe63d[1][1]} + {irbe63d[1][2][ym3b97e-1],irbe63d[1][2]};               aabc866[1] <=  {qt6f1bc[1][vk2fc20-1],qt6f1bc[1]}     + {wjc6f21[1][vk2fc20-1],wjc6f21[1]};
               qt6f1bc[2] <=  ui56a8c;               wjc6f21[2] <=  {irbe63d[2][1][ym3b97e-1],irbe63d[2][1]} + {irbe63d[2][2][ym3b97e-1],irbe63d[2][2]};               aabc866[2] <=  {qt6f1bc[2][vk2fc20-1],qt6f1bc[2]}     + {wjc6f21[2][vk2fc20-1],wjc6f21[2]};            end         end      end   end else if (CORETYPE == 13) begin        always @(posedge clk or negedge rstn) begin         if (!rstn) begin            aabc866[0] <= {gof081f{1'b0}} ;            aabc866[1] <= {gof081f{1'b0}} ;            aabc866[2] <= {gof081f{1'b0}} ;         end else if (ngb77c) begin            if (kd5bbe3) begin               aabc866[0] <= {gof081f{1'b0}} ;               aabc866[1] <= {gof081f{1'b0}} ;               aabc866[2] <= {gof081f{1'b0}} ;            end else begin               aabc866[0] <=  {ui56a8c[vk2fc20-1],ui56a8c};               aabc866[1] <=  {irbe63d[1][1][ym3b97e-1],irbe63d[1][1][ym3b97e-1],irbe63d[1][1]} +                               {irbe63d[1][2][ym3b97e-1],irbe63d[1][2][ym3b97e-1],irbe63d[1][2]};               aabc866[2] <=  {irbe63d[2][1][ym3b97e-1],irbe63d[2][1][ym3b97e-1],irbe63d[2][1]} +                               {irbe63d[2][2][ym3b97e-1],irbe63d[2][2][ym3b97e-1],irbe63d[2][2]};            end         end      end   end
end
endgenerate
assign dout0 = aabc866[0];
assign dout1 = aabc866[1];
assign dout2 = aabc866[2];
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];jc7c771<={din0>>1,fp2dc72[2]};oh1dc57<={din1>>1,fp2dc72[3]};jp715e2<={din2>>1,fp2dc72[4]};ui56a8c<={ou98f6f>>1,fp2dc72[5]};xlaa30e<={ym2198b>>1,fp2dc72[6]};tw8c3b4<={ho662c7>>1,fp2dc72[7]};pued16<={fp8b1d0>>1,fp2dc72[8]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=din0[0];vk25b8e[2044]<=din1[0];vk25b8e[2041]<=din2[0];vk25b8e[2035]<=ou98f6f[0];vk25b8e[2022]<=ym2198b[0];vk25b8e[1996]<=ho662c7[0];vk25b8e[1945]<=fp8b1d0[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module rv6684_colorspace (
                     clk,   
                     rstn,
                     ce,
                     sr,
                     din0,
                     din1,
                     din2,
                     dout0,
                     dout1,
                     dout2);
parameter      CORETYPE          = 0;
parameter      psdaa9a        = 12;
parameter      CWIDTH            = 8;
parameter      CPOINTS           = 0;
parameter      ym3b97e      = 20;
parameter      vk2fc20    = 21;
parameter      gof081f    = 22;
parameter      DINSIGN           = "Signed";
parameter      DSPBLKMULT        = "Enable";
parameter      INSERIAL          = "Serial";
parameter      DEVICE            = "ECP2";
parameter      CV_MH             = 0;
parameter      CV_MI             = 0;
parameter      CV_MJ             = 0;
parameter      CV_MK             = 0;
parameter      CV_NH             = 0;
parameter      CV_NI             = 0;
parameter      CV_NJ             = 0;
parameter      CV_NK             = 0;
parameter      CV_PH             = 0;
parameter      CV_PI             = 0;
parameter      CV_PJ             = 0;
parameter      CV_PK             = 0;
localparam     fae46b8    = (DINSIGN == "Signed")? (psdaa9a+1) : (psdaa9a+2);
localparam     ngb870e      = fae46b8;
localparam     jr1c394      = ngb870e + CWIDTH;
localparam     qg729d3      = jr1c394 + 1;
localparam     baa74c6      = qg729d3 + 1;
localparam     ald3193      = gof081f - CWIDTH ;
input                               clk;
input                               rstn;
input                               ce;
input                               sr;
input        [psdaa9a-1:0]       din0;
input        [psdaa9a-1:0]       din1;
input        [psdaa9a-1:0]       din2;
output       [gof081f-1:0]   dout0;
output       [gof081f-1:0]   dout1;
output       [gof081f-1:0]   dout2;
wire         [CWIDTH-1:0]           th5ae22 [0:2][0:2];
wire         [fae46b8-1:0]   tufe57d;
wire         [fae46b8-1:0]   gd95f5c;
wire         [fae46b8-1:0]   cm7d727;
wire         [fae46b8-1:0]   fp8b1d0;
wire         [fae46b8-1:0]   zz270c2;
wire         [fae46b8-1:0]   ofc30b6;
wire                                oh185b5;
wire                                blc2dad;
wire         [gof081f-2:0]   wyb6b77;
wire         [gof081f-2:0]   puaddc7;
wire         [gof081f-1:0]   yk771d7;
wire         [gof081f-1:0]   jpc75cb;
wire         [gof081f-1:0]   xjd72fa;
wire                                ksb97d6;
wire                                eacbeb0;
wire         [psdaa9a-1:0]       mefac06;
wire         [psdaa9a-1:0]       fpb0184;
wire         [psdaa9a:0]         ph6135;
wire         [psdaa9a:0]         rv84d7b;
wire         [psdaa9a:0]         ng35efd;
wire         [jr1c394-1:0]     ld7bf5e;
wire         [jr1c394-1:0]     shfd7b3;
wire         [gof081f-1:0]   gb5ece3;
wire         [gof081f-1:0]   swb38ef;
wire         [jr1c394-1:0]     the3bc3;
wire         [jr1c394-1:0]     ayef0fc;
wire         [gof081f-1:0]   dout0;
wire         [gof081f-1:0]   dout1;
wire         [gof081f-1:0]   dout2;
reg          [psdaa9a-1:0]       ou98f6f[0:5];
reg          [psdaa9a-1:0]       pf71283[0:5];
reg          [psdaa9a-1:0]       xj4a0f2[0:5];
reg          [ngb870e-1:0]     ng83cbf;
reg          [ngb870e-1:0]     wjf2fd2;
reg          [ngb870e-1:0]     dbbf4a1;
reg          [ngb870e-1:0]     pfd2879;
reg          [qg729d3-1:0]     cba1e7f;
reg          [baa74c6-1:0]     fa79fe1;
reg          [ald3193-1:0]     sh7f85a;
reg          [ald3193-1:0]     zke16a6;
reg          [ald3193-1:0]     ld5a99b;
reg          [ald3193-1:0]     iea66f8;
reg          [gof081f-1:0]   lf9be05;
reg          [gof081f-1:0]   wjf817a;
reg          [gof081f-1:0]   gq5ea3;
reg          [gof081f-1:0]   en7a8ca;
reg          [jr1c394-1:0]     yma32a1;
reg          [jr1c394-1:0]     psca847;
reg          [gof081f-1:0]   ira11d5;
reg          [gof081f-1:0]   vi4756d;
integer cm4915d;
reg ngb77c;
reg kd5bbe3;
reg [psdaa9a - 1 : 0] jc7c771;
reg [psdaa9a - 1 : 0] oh1dc57;
reg [psdaa9a - 1 : 0] jp715e2;
reg [fae46b8 - 1 : 0] ho76c36;
reg [fae46b8 - 1 : 0] vxb0d91;
reg [fae46b8 - 1 : 0] sj3647a;
reg [fae46b8 - 1 : 0] pued16;
reg [fae46b8 - 1 : 0] of7aaf5;
reg [fae46b8 - 1 : 0] yzabd63;
reg kd5eb1d;
reg suf58ed;
reg [gof081f - 2 : 0] xw63b49;
reg [gof081f - 2 : 0] yxed25c;
reg [gof081f - 1 : 0] su4972b;
reg [gof081f - 1 : 0] ic5cac4;
reg [gof081f - 1 : 0] ec2b101;
reg by58808;
reg uic4042;
reg [psdaa9a - 1 : 0] je1083;
reg [psdaa9a - 1 : 0] zk420d4;
reg [psdaa9a : 0] hq83519;
reg [psdaa9a : 0] cmd4659;
reg [psdaa9a : 0] jr19648;
reg [jr1c394 - 1 : 0] kq59239;
reg [jr1c394 - 1 : 0] jc48e4c;
reg [gof081f - 1 : 0] ep3931b;
reg [gof081f - 1 : 0] kq4c6e5;
reg [jr1c394 - 1 : 0] vk1b942;
reg [jr1c394 - 1 : 0] sue509c;
reg [ngb870e - 1 : 0] jc4270f;
reg [ngb870e - 1 : 0] vk9c3df;
reg [ngb870e - 1 : 0] ouf7da;
reg [ngb870e - 1 : 0] zkdf68e;
reg [qg729d3 - 1 : 0] vida393;
reg [baa74c6 - 1 : 0] vx8e4d0;
reg [ald3193 - 1 : 0] hq93439;
reg [ald3193 - 1 : 0] vid0e54;
reg [ald3193 - 1 : 0] kf39511;
reg [ald3193 - 1 : 0] uv54462;
reg [gof081f - 1 : 0] xy118aa;
reg [gof081f - 1 : 0] os62a92;
reg [gof081f - 1 : 0] fpaa489;
reg [gof081f - 1 : 0] co92272;
reg [jr1c394 - 1 : 0] vk89c87;
reg [jr1c394 - 1 : 0] cm721dd;
reg [gof081f - 1 : 0] mg8774c;
reg [gof081f - 1 : 0] zxdd308;
reg [2047:0] vk25b8e;
wire [48:0] fp2dc72;
localparam ld6e396 = 49,hb71cb6 = 32'hfdffd84b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
assign       th5ae22[0][0] = CV_MH ;
assign       th5ae22[0][1] = CV_MI ;
assign       th5ae22[0][2] = CV_MJ ;
assign       th5ae22[1][0] = CV_NH ;
assign       th5ae22[1][1] = CV_NI ;
assign       th5ae22[1][2] = CV_NJ ;
assign       th5ae22[2][0] = CV_PH ;
assign       th5ae22[2][1] = CV_PI ;
assign       th5ae22[2][2] = CV_PJ ;
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      for (cm4915d=0;cm4915d<6;cm4915d=cm4915d+1) begin : ep887a         ou98f6f[cm4915d] <= {psdaa9a{1'b0}};         pf71283[cm4915d] <= {psdaa9a{1'b0}};         xj4a0f2[cm4915d] <= {psdaa9a{1'b0}};      end   end else if (ngb77c) begin      if (kd5bbe3) begin         for (cm4915d=0;cm4915d<6;cm4915d=cm4915d+1) begin : ec821e0            ou98f6f[cm4915d] <= {psdaa9a{1'b0}};            pf71283[cm4915d] <= {psdaa9a{1'b0}};            xj4a0f2[cm4915d] <= {psdaa9a{1'b0}};         end      end else begin         ou98f6f[0] <= jc7c771;         pf71283[0] <= oh1dc57;         xj4a0f2[0] <= jp715e2;         for (cm4915d=1;cm4915d<6;cm4915d=cm4915d+1) begin : mrc99b3            ou98f6f[cm4915d] <= ou98f6f[cm4915d-1];            pf71283[cm4915d] <= pf71283[cm4915d-1];            xj4a0f2[cm4915d] <= xj4a0f2[cm4915d-1];         end      end   end
end
assign tufe57d = (DINSIGN == "Signed") ? {jc7c771[psdaa9a-1],jc7c771} : {2'b00,jc7c771};
assign gd95f5c = (DINSIGN == "Signed") ? {oh1dc57[psdaa9a-1],oh1dc57} : {2'b00,oh1dc57};
assign cm7d727 = (DINSIGN == "Signed") ? {jp715e2[psdaa9a-1],jp715e2} : {2'b00,jp715e2};
assign fp8b1d0  = (DINSIGN == "Signed") ? {ou98f6f[5][psdaa9a-1],ou98f6f[5]} : {2'b00,ou98f6f[5]};
assign zz270c2  = (DINSIGN == "Signed") ? {pf71283[4][psdaa9a-1],pf71283[4]} : {2'b00,pf71283[4]};
assign ofc30b6  = (DINSIGN == "Signed") ? {xj4a0f2[5][psdaa9a-1],xj4a0f2[5]} : {2'b00,xj4a0f2[5]};
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      ng83cbf  <=  {ngb870e{1'b0}};      wjf2fd2 <=  {ngb870e{1'b0}};      dbbf4a1  <=  {ngb870e{1'b0}};      pfd2879 <=  {ngb870e{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         ng83cbf  <=  {ngb870e{1'b0}};         wjf2fd2 <=  {ngb870e{1'b0}};         dbbf4a1  <=  {ngb870e{1'b0}};         pfd2879 <=  {ngb870e{1'b0}};      end else begin         ng83cbf  <=  ho76c36 - vxb0d91;         wjf2fd2 <=  jc4270f;         dbbf4a1  <=  sj3647a - vxb0d91;         pfd2879 <=  ouf7da;      end   end
end
generate begin   if (DSPBLKMULT == "Enable") begin       pmi_dsp_mult   #(.pmi_dataa_width           (ngb870e   ),                        .pmi_datab_width           (CWIDTH         ),                        .pmi_additional_pipeline   (1              ),                        .pmi_input_reg             ("on"           ),                        .pmi_output_reg            ("on"           ),                        .pmi_family                (DEVICE         ),                        .pmi_gsr                   ("enable"       ),                        .pmi_source_control_a      ("parallel"     ),                        .pmi_source_control_b      ("parallel"     ),                        .pmi_reg_inputa_clk        ("CLK0"         ),                        .pmi_reg_inputa_ce         ("CE0"          ),                        .pmi_reg_inputa_rst        ("RST0"         ),                        .pmi_reg_inputb_clk        ("CLK0"         ),                        .pmi_reg_inputb_ce         ("CE0"          ),                        .pmi_reg_inputb_rst        ("RST0"         ),                        .pmi_reg_pipeline_clk      ("CLK0"         ),                        .pmi_reg_pipeline_ce       ("CE0"          ),                        .pmi_reg_pipeline_rst      ("RST0"         ),                        .pmi_reg_output_clk        ("CLK0"         ),                        .pmi_reg_output_ce         ("CE0"          ),                        .pmi_reg_output_rst        ("RST0"         ),                        .pmi_reg_signeda_clk       ("CLK0"         ),                        .pmi_reg_signeda_ce        ("CE0"          ),                        .pmi_reg_signeda_rst       ("RST0"         ),                        .pmi_reg_signedb_clk       ("CLK0"         ),                        .pmi_reg_signedb_ce        ("CE0"          ),                        .pmi_reg_signedb_rst       ("RST0"         ),                        .pmi_pipelined_mode        ("off"          ),                        .module_type               ("pmi_dsp_mult" ))       zx5565d  (                        .A                         (ng83cbf         ),                        .B                         (th5ae22[0][1]       ),                        .SRIA                      (               ),                        .SRIB                      (               ),                        .CLK0                      (clk            ),                        .CLK1                      (clk            ),                        .CLK2                      (clk            ),                        .CLK3                      (clk            ),                        .CE0                       (ce             ),                        .CE1                       (ce             ),                        .CE2                       (ce             ),                        .CE3                       (ce             ),                        .RST0                      (~rstn          ),                        .RST1                      (~rstn          ),                        .RST2                      (~rstn          ),                        .RST3                      (~rstn          ),                        .SignA                     (1'b1           ),                        .SignB                     (1'b1           ),                        .SourceA                   (1'b0           ),                        .SourceB                   (1'b0           ),                        .P                         (the3bc3   ),                        .SROA                      (               ),                        .SROB                      (               ));       pmi_dsp_mult   #(.pmi_dataa_width           (ngb870e   ),                        .pmi_datab_width           (CWIDTH         ),                        .pmi_additional_pipeline   (1              ),                        .pmi_input_reg             ("on"           ),                        .pmi_output_reg            ("on"           ),                        .pmi_family                (DEVICE         ),                        .pmi_gsr                   ("enable"       ),                        .pmi_source_control_a      ("parallel"     ),                        .pmi_source_control_b      ("parallel"     ),                        .pmi_reg_inputa_clk        ("CLK0"         ),                        .pmi_reg_inputa_ce         ("CE0"          ),                        .pmi_reg_inputa_rst        ("RST0"         ),                        .pmi_reg_inputb_clk        ("CLK0"         ),                        .pmi_reg_inputb_ce         ("CE0"          ),                        .pmi_reg_inputb_rst        ("RST0"         ),                        .pmi_reg_pipeline_clk      ("CLK0"         ),                        .pmi_reg_pipeline_ce       ("CE0"          ),                        .pmi_reg_pipeline_rst      ("RST0"         ),                        .pmi_reg_output_clk        ("CLK0"         ),                        .pmi_reg_output_ce         ("CE0"          ),                        .pmi_reg_output_rst        ("RST0"         ),                        .pmi_reg_signeda_clk       ("CLK0"         ),                        .pmi_reg_signeda_ce        ("CE0"          ),                        .pmi_reg_signeda_rst       ("RST0"         ),                        .pmi_reg_signedb_clk       ("CLK0"         ),                        .pmi_reg_signedb_ce        ("CE0"          ),                        .pmi_reg_signedb_rst       ("RST0"         ),                        .pmi_pipelined_mode        ("off"          ),                        .module_type               ("pmi_dsp_mult" ))       en5e7fc  (                        .A                         (dbbf4a1         ),                        .B                         (th5ae22[0][2]       ),                        .SRIA                      (               ),                        .SRIB                      (               ),                        .CLK0                      (clk            ),                        .CLK1                      (clk            ),                        .CLK2                      (clk            ),                        .CLK3                      (clk            ),                        .CE0                       (ce             ),                        .CE1                       (ce             ),                        .CE2                       (ce             ),                        .CE3                       (ce             ),                        .RST0                      (~rstn          ),                        .RST1                      (~rstn          ),                        .RST2                      (~rstn          ),                        .RST3                      (~rstn          ),                        .SignA                     (1'b1           ),                        .SignB                     (1'b1           ),                        .SourceA                   (1'b0           ),                        .SourceB                   (1'b0           ),                        .P                         (ayef0fc   ),                        .SROA                      (               ),                        .SROB                      (               ));
       pmi_dsp_mult   #(.pmi_dataa_width           (ald3193   ),                        .pmi_datab_width           (CWIDTH         ),                        .pmi_additional_pipeline   (1              ),                        .pmi_input_reg             ("on"           ),                        .pmi_output_reg            ("on"           ),                        .pmi_family                (DEVICE         ),                        .pmi_gsr                   ("enable"       ),                        .pmi_source_control_a      ("parallel"     ),                        .pmi_source_control_b      ("parallel"     ),                        .pmi_reg_inputa_clk        ("CLK0"         ),                        .pmi_reg_inputa_ce         ("CE0"          ),                        .pmi_reg_inputa_rst        ("RST0"         ),                        .pmi_reg_inputb_clk        ("CLK0"         ),                        .pmi_reg_inputb_ce         ("CE0"          ),                        .pmi_reg_inputb_rst        ("RST0"         ),                        .pmi_reg_pipeline_clk      ("CLK0"         ),                        .pmi_reg_pipeline_ce       ("CE0"          ),                        .pmi_reg_pipeline_rst      ("RST0"         ),                        .pmi_reg_output_clk        ("CLK0"         ),                        .pmi_reg_output_ce         ("CE0"          ),                        .pmi_reg_output_rst        ("RST0"         ),                        .pmi_reg_signeda_clk       ("CLK0"         ),                        .pmi_reg_signeda_ce        ("CE0"          ),                        .pmi_reg_signeda_rst       ("RST0"         ),                        .pmi_reg_signedb_clk       ("CLK0"         ),                        .pmi_reg_signedb_ce        ("CE0"          ),                        .pmi_reg_signedb_rst       ("RST0"         ),                        .pmi_pipelined_mode        ("off"          ),                        .module_type               ("pmi_dsp_mult" ))       gq92975  (                        .A                         (sh7f85a         ),                        .B                         (th5ae22[1][0]       ),                        .SRIA                      (               ),                        .SRIB                      (               ),                        .CLK0                      (clk            ),                        .CLK1                      (clk            ),                        .CLK2                      (clk            ),                        .CLK3                      (clk            ),                        .CE0                       (ce             ),                        .CE1                       (ce             ),                        .CE2                       (ce             ),                        .CE3                       (ce             ),                        .RST0                      (~rstn          ),                        .RST1                      (~rstn          ),                        .RST2                      (~rstn          ),                        .RST3                      (~rstn          ),                        .SignA                     (1'b1           ),                        .SignB                     (1'b1           ),                        .SourceA                   (1'b0           ),                        .SourceB                   (1'b0           ),                        .P                         (dout1          ),                        .SROA                      (               ),                        .SROB                      (               ));       pmi_dsp_mult   #(.pmi_dataa_width           (ald3193   ),                        .pmi_datab_width           (CWIDTH         ),                        .pmi_additional_pipeline   (1              ),                        .pmi_input_reg             ("on"           ),                        .pmi_output_reg            ("on"           ),                        .pmi_family                (DEVICE         ),                        .pmi_gsr                   ("enable"       ),                        .pmi_source_control_a      ("parallel"     ),                        .pmi_source_control_b      ("parallel"     ),                        .pmi_reg_inputa_clk        ("CLK0"         ),                        .pmi_reg_inputa_ce         ("CE0"          ),                        .pmi_reg_inputa_rst        ("RST0"         ),                        .pmi_reg_inputb_clk        ("CLK0"         ),                        .pmi_reg_inputb_ce         ("CE0"          ),                        .pmi_reg_inputb_rst        ("RST0"         ),                        .pmi_reg_pipeline_clk      ("CLK0"         ),                        .pmi_reg_pipeline_ce       ("CE0"          ),                        .pmi_reg_pipeline_rst      ("RST0"         ),                        .pmi_reg_output_clk        ("CLK0"         ),                        .pmi_reg_output_ce         ("CE0"          ),                        .pmi_reg_output_rst        ("RST0"         ),                        .pmi_reg_signeda_clk       ("CLK0"         ),                        .pmi_reg_signeda_ce        ("CE0"          ),                        .pmi_reg_signeda_rst       ("RST0"         ),                        .pmi_reg_signedb_clk       ("CLK0"         ),                        .pmi_reg_signedb_ce        ("CE0"          ),                        .pmi_reg_signedb_rst       ("RST0"         ),                        .pmi_pipelined_mode        ("off"          ),                        .module_type               ("pmi_dsp_mult" ))       fa69ac3  (                        .A                         (ld5a99b         ),                        .B                         (th5ae22[2][0]       ),                        .SRIA                      (               ),                        .SRIB                      (               ),                        .CLK0                      (clk            ),                        .CLK1                      (clk            ),                        .CLK2                      (clk            ),                        .CLK3                      (clk            ),                        .CE0                       (ce             ),                        .CE1                       (ce             ),                        .CE2                       (ce             ),                        .CE3                       (ce             ),                        .RST0                      (~rstn          ),                        .RST1                      (~rstn          ),                        .RST2                      (~rstn          ),                        .RST3                      (~rstn          ),                        .SignA                     (1'b1           ),                        .SignB                     (1'b1           ),                        .SourceA                   (1'b0           ),                        .SourceB                   (1'b0           ),                        .P                         (dout2          ),                        .SROA                      (               ),                        .SROB                      (               ));   end else begin                     always @(posedge clk or negedge rstn) begin                        if (!rstn) begin                           yma32a1 <= {jr1c394{1'b0}};                        end else if (ngb77c) begin                           if (kd5bbe3) begin                              yma32a1 <= {jr1c394{1'b0}};                           end else begin                              yma32a1 <= kq59239;                           end                         end                     end                     db199ce_colorspace # (.psdaa9a                (ngb870e        ),                              .sj39da8                 (CWIDTH              ),                              .jc76a28                     ("Signed"            ),                              .lsa8a16                     ("Signed"            ))                    qv12a54 (.clk                       (clk                 ),                              .rstn                      (rstn                ),
                              .ce                        (ngb77c                  ),                              .sr                        (kd5bbe3                  ),                              .pub26f4                  (jc4270f              ),                              .uide8d7                  (th5ae22[0][1]            ),                              .irbe63d                  (ld7bf5e          ));
                     assign the3bc3 = vk89c87;
                     always @(posedge clk or negedge rstn) begin                        if (!rstn) begin                           psca847 <= {jr1c394{1'b0}};                        end else if (ngb77c) begin                           if (kd5bbe3) begin                              psca847 <= {jr1c394{1'b0}};                           end else begin                              psca847 <= jc48e4c;                           end                         end                     end                     db199ce_colorspace # (.psdaa9a                (ngb870e        ),                              .sj39da8                 (CWIDTH              ),                              .jc76a28                     ("Signed"            ),                              .lsa8a16                     ("Signed"            ))                    uk825f4 (.clk                       (clk                 ),                              .rstn                      (rstn                ),                              .ce                        (ngb77c                  ),                              .sr                        (kd5bbe3                  ),                              .pub26f4                  (ouf7da              ),                              .uide8d7                  (th5ae22[0][2]            ),                              .irbe63d                  (shfd7b3          ));
                     assign ayef0fc = cm721dd;
                     always @(posedge clk or negedge rstn) begin                        if (!rstn) begin                           ira11d5 <= {gof081f{1'b0}};                        end else if (ngb77c) begin                           if (kd5bbe3) begin                              ira11d5 <= {gof081f{1'b0}};                           end else begin                              ira11d5 <= ep3931b;                           end                         end                     end                     db199ce_colorspace # (.psdaa9a                (ald3193        ),                              .sj39da8                 (CWIDTH              ),                              .jc76a28                     ("Signed"            ),                              .lsa8a16                     ("Signed"            ))                    vvf9c5d (.clk                       (clk                 ),                              .rstn                      (rstn                ),                              .ce                        (ngb77c                  ),                              .sr                        (kd5bbe3                  ),                              .pub26f4                  (hq93439              ),                              .uide8d7                  (th5ae22[1][0]            ),                              .irbe63d                  (gb5ece3          ));
                     assign dout1 = mg8774c;                     always @(posedge clk or negedge rstn) begin                        if (!rstn) begin                           vi4756d <= {gof081f{1'b0}};                        end else if (ngb77c) begin                           if (kd5bbe3) begin                              vi4756d <= {gof081f{1'b0}};                           end else begin                              vi4756d <= kq4c6e5;                           end                         end                     end                     db199ce_colorspace # (.psdaa9a                (ald3193        ),                              .sj39da8                 (CWIDTH              ),                              .jc76a28                     ("Signed"            ),                              .lsa8a16                     ("Signed"            ))                    hofe0f5 (.clk                       (clk                 ),                              .rstn                      (rstn                ),                              .ce                        (ngb77c                  ),                              .sr                        (kd5bbe3                  ),                              .pub26f4                  (kf39511              ),                              .uide8d7                  (th5ae22[2][0]            ),                              .irbe63d                  (swb38ef          ));
                     assign dout2 = zxdd308;
   end      always @(posedge clk or negedge rstn) begin         if (!rstn) begin            sh7f85a  <= {ald3193{1'b0}};            zke16a6 <= {ald3193{1'b0}};            ld5a99b  <= {ald3193{1'b0}};            iea66f8 <= {ald3193{1'b0}};         end else if (ngb77c) begin            if (kd5bbe3) begin               sh7f85a  <= {ald3193{1'b0}};               zke16a6 <= {ald3193{1'b0}};               ld5a99b  <= {ald3193{1'b0}};               iea66f8 <= {ald3193{1'b0}};            end else begin               if (ald3193 == fae46b8) begin                  sh7f85a  <= yzabd63 - {jr19648[psdaa9a],jr19648};                  zke16a6 <= hq93439;                  ld5a99b  <= pued16 - {jr19648[psdaa9a],jr19648};                  iea66f8 <= kf39511;               end else begin                  sh7f85a  <=  {{(ald3193-fae46b8){yzabd63[fae46b8-1]}},yzabd63} - {jr19648[psdaa9a],jr19648};                  zke16a6 <= hq93439;                  ld5a99b  <= {{(ald3193-fae46b8){pued16[fae46b8-1]}},pued16} - {jr19648[psdaa9a],jr19648};                  iea66f8 <= kf39511;               end            end         end      end
end
endgenerate
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      cba1e7f <=  {qg729d3{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         cba1e7f <=  {qg729d3{1'b0}};      end else begin         cba1e7f <=  {vk1b942[jr1c394-1],vk1b942} + {sue509c[jr1c394-1],sue509c} ;      end   end
end
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      fa79fe1 <=  {baa74c6{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         fa79fe1 <=  {baa74c6{1'b0}};      end else begin         fa79fe1 <= {vida393[qg729d3-1],vida393} + {{(baa74c6-fae46b8-CPOINTS){of7aaf5[fae46b8-1]}},of7aaf5,{CPOINTS{1'b0}}};      end   end
end
assign wyb6b77    = {(gof081f-1){1'b0}};
assign puaddc7     = {(gof081f-1){1'b1}};
assign oh185b5  = |(vx8e4d0[baa74c6-1:gof081f-1]);
assign blc2dad = &(vx8e4d0[baa74c6-1:gof081f-1]);
assign yk771d7    = suf58ed ? vx8e4d0[gof081f-1:0] : {1'b1,xw63b49};
assign jpc75cb    = kd5eb1d ? {1'b0,yxed25c} : vx8e4d0[gof081f-1:0];
assign xjd72fa    = vx8e4d0[baa74c6-1] ? su4972b : ic5cac4;
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      lf9be05 <= {gof081f{1'b0}};      wjf817a <= {gof081f{1'b0}};      gq5ea3 <= {gof081f{1'b0}};      en7a8ca <= {gof081f{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         lf9be05 <= {gof081f{1'b0}};         wjf817a <= {gof081f{1'b0}};         gq5ea3 <= {gof081f{1'b0}};         en7a8ca <= {gof081f{1'b0}};      end else begin         lf9be05 <= ec2b101;         wjf817a <= xy118aa;         gq5ea3 <= os62a92;         en7a8ca <= fpaa489;      end   end
end
assign dout0 = co92272;
assign mefac06    = {psdaa9a{1'b0}};
assign fpb0184     = {psdaa9a{1'b1}};
assign ksb97d6  = |(vx8e4d0[baa74c6-1:psdaa9a+CPOINTS]);
assign eacbeb0 = &(vx8e4d0[baa74c6-1:psdaa9a+CPOINTS]);
assign ph6135    = uic4042 ? vx8e4d0[psdaa9a+CPOINTS:CPOINTS] : {1'b1,je1083};
assign rv84d7b    = by58808 ? {1'b0,zk420d4} : vx8e4d0[psdaa9a+CPOINTS:CPOINTS];
assign ng35efd    = vx8e4d0[baa74c6-1] ? hq83519 : cmd4659;
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];jc7c771<={din0>>1,fp2dc72[2]};oh1dc57<={din1>>1,fp2dc72[3]};jp715e2<={din2>>1,fp2dc72[4]};ho76c36<={tufe57d>>1,fp2dc72[5]};vxb0d91<={gd95f5c>>1,fp2dc72[6]};sj3647a<={cm7d727>>1,fp2dc72[7]};pued16<={fp8b1d0>>1,fp2dc72[8]};of7aaf5<={zz270c2>>1,fp2dc72[9]};yzabd63<={ofc30b6>>1,fp2dc72[10]};kd5eb1d<=fp2dc72[11];suf58ed<=fp2dc72[12];xw63b49<={wyb6b77>>1,fp2dc72[13]};yxed25c<={puaddc7>>1,fp2dc72[14]};su4972b<={yk771d7>>1,fp2dc72[15]};ic5cac4<={jpc75cb>>1,fp2dc72[16]};ec2b101<={xjd72fa>>1,fp2dc72[17]};by58808<=fp2dc72[18];uic4042<=fp2dc72[19];je1083<={mefac06>>1,fp2dc72[20]};zk420d4<={fpb0184>>1,fp2dc72[21]};hq83519<={ph6135>>1,fp2dc72[22]};cmd4659<={rv84d7b>>1,fp2dc72[23]};jr19648<={ng35efd>>1,fp2dc72[24]};kq59239<={ld7bf5e>>1,fp2dc72[25]};jc48e4c<={shfd7b3>>1,fp2dc72[26]};ep3931b<={gb5ece3>>1,fp2dc72[27]};kq4c6e5<={swb38ef>>1,fp2dc72[28]};vk1b942<={the3bc3>>1,fp2dc72[29]};sue509c<={ayef0fc>>1,fp2dc72[30]};jc4270f<={ng83cbf>>1,fp2dc72[31]};vk9c3df<={wjf2fd2>>1,fp2dc72[32]};ouf7da<={dbbf4a1>>1,fp2dc72[33]};zkdf68e<={pfd2879>>1,fp2dc72[34]};vida393<={cba1e7f>>1,fp2dc72[35]};vx8e4d0<={fa79fe1>>1,fp2dc72[36]};hq93439<={sh7f85a>>1,fp2dc72[37]};vid0e54<={zke16a6>>1,fp2dc72[38]};kf39511<={ld5a99b>>1,fp2dc72[39]};uv54462<={iea66f8>>1,fp2dc72[40]};xy118aa<={lf9be05>>1,fp2dc72[41]};os62a92<={wjf817a>>1,fp2dc72[42]};fpaa489<={gq5ea3>>1,fp2dc72[43]};co92272<={en7a8ca>>1,fp2dc72[44]};vk89c87<={yma32a1>>1,fp2dc72[45]};cm721dd<={psca847>>1,fp2dc72[46]};mg8774c<={ira11d5>>1,fp2dc72[47]};zxdd308<={vi4756d>>1,fp2dc72[48]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=din0[0];vk25b8e[2044]<=din1[0];vk25b8e[2040]<=din2[0];vk25b8e[2033]<=tufe57d[0];vk25b8e[2019]<=gd95f5c[0];vk25b8e[1999]<=cba1e7f[0];vk25b8e[1991]<=cm7d727[0];vk25b8e[1950]<=fa79fe1[0];vk25b8e[1947]<=wjf817a[0];vk25b8e[1934]<=fp8b1d0[0];vk25b8e[1892]<=mefac06[0];vk25b8e[1852]<=sh7f85a[0];vk25b8e[1851]<=yk771d7[0];vk25b8e[1847]<=gq5ea3[0];vk25b8e[1820]<=zz270c2[0];vk25b8e[1783]<=vi4756d[0];vk25b8e[1737]<=fpb0184[0];vk25b8e[1657]<=zke16a6[0];vk25b8e[1654]<=jpc75cb[0];vk25b8e[1647]<=en7a8ca[0];vk25b8e[1610]<=ng35efd[0];vk25b8e[1593]<=ofc30b6[0];vk25b8e[1523]<=dbbf4a1[0];vk25b8e[1426]<=ph6135[0];vk25b8e[1404]<=ng83cbf[0];vk25b8e[1267]<=ld5a99b[0];vk25b8e[1260]<=xjd72fa[0];vk25b8e[1246]<=yma32a1[0];vk25b8e[1199]<=swb38ef[0];vk25b8e[1173]<=ld7bf5e[0];vk25b8e[1139]<=oh185b5;vk25b8e[1023]<=ce;vk25b8e[999]<=pfd2879[0];vk25b8e[973]<=lf9be05[0];vk25b8e[946]<=eacbeb0;vk25b8e[925]<=puaddc7[0];vk25b8e[891]<=ira11d5[0];vk25b8e[805]<=rv84d7b[0];vk25b8e[761]<=wjf2fd2[0];vk25b8e[702]<=ayef0fc[0];vk25b8e[599]<=gb5ece3[0];vk25b8e[486]<=iea66f8[0];vk25b8e[473]<=ksb97d6;vk25b8e[462]<=wyb6b77[0];vk25b8e[445]<=psca847[0];vk25b8e[351]<=the3bc3[0];vk25b8e[299]<=shfd7b3[0];vk25b8e[231]<=blc2dad;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module xy1b553_colorspace (
               
               clk,                 
               rstn,                
               ce,                  
               sr,                  
               ph27078,                 
               
               wwc1e36                 
               );
parameter psdaa9a             =8;
input                                     clk;
input                                     rstn;
input                                     ce;
input                                     sr;
input  [psdaa9a-1:0]                   ph27078;
output [psdaa9a-1:0]                   wwc1e36;
reg    [psdaa9a-1:0]                   wwc1e36;
reg ngb77c;
reg kd5bbe3;
reg [psdaa9a - 1 : 0] wy15935;
reg [2047:0] vk25b8e;
wire [2:0] fp2dc72;
localparam ld6e396 = 3,hb71cb6 = 32'hfdffc70b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
always @(posedge clk or negedge rstn) begin   if (!rstn)      wwc1e36 <= 0;   else if (ngb77c) begin      if (kd5bbe3)         wwc1e36 <= {psdaa9a{1'b0}};      else         wwc1e36 <= wy15935;   end
end
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];wy15935<={ph27078>>1,fp2dc72[2]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=ph27078[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module twa8e69_colorspace (
             
             clk,
             rstn,
             ce,
             sr,
             ph27078,
             
             wwc1e36
             );
parameter yz39132           = 12;
parameter DOUTWIDTH        = 32;
parameter sw212c2    = 1;
parameter ph329ec    = "Rounding away from zero";
parameter al44ca7    = "Saturation";
parameter yx70b70            = 24;
parameter ps66cfe        = 0;
parameter CPOINTS          = 0;
parameter DOUTPOINTS       = 0;
parameter pua7b36         = "Signed";
parameter nt3d9b3        = "Signed";
parameter ene8af1         = 0;
localparam uxabeb4 = (DOUTPOINTS < ps66cfe+CPOINTS) ? ps66cfe+CPOINTS-DOUTPOINTS : 0;
localparam eaea539 = (uxabeb4 == 0) ? yz39132 :                       (ph329ec == "Truncation") ? yz39132-uxabeb4 :                       (pua7b36 == "Unsigned") ? yz39132-uxabeb4+1 : yz39132-uxabeb4+2;
localparam gq92cf6 = (DOUTPOINTS>=(ps66cfe+CPOINTS)) ? (DOUTWIDTH+ps66cfe+CPOINTS-DOUTPOINTS) :                        ((DOUTWIDTH>(yz39132-uxabeb4)) ? (yz39132-uxabeb4) : DOUTWIDTH);
localparam oh85b85 = (pua7b36 == "Unsigned") ? yz39132-uxabeb4 : yz39132-uxabeb4+1;
localparam dz6ed6e = (oh85b85+yx70b70-1)/yx70b70;
input                       clk;
input                       rstn;
input                       ce;
input                       sr;
input[yz39132-1:0]           ph27078;
output [DOUTWIDTH-1:0]      wwc1e36;
wire[eaea539-1:0]         tj9ee2b;
reg[yz39132-1:0]             lsb8afd;
reg ngb77c;
reg kd5bbe3;
reg [yz39132 - 1 : 0] wy15935;
reg [eaea539 - 1 : 0] bl5a3e2;
reg [yz39132 - 1 : 0] oh8f8b0;
reg [2047:0] vk25b8e;
wire [4:0] fp2dc72;
localparam ld6e396 = 5,hb71cb6 = 32'hfdffe0cb;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
generate
begin   if (ene8af1 == 1) begin      always @(posedge clk or negedge rstn)      begin         if (rstn == 1'b0)            lsb8afd <= {yz39132{1'b0}};         else if (ngb77c == 1'b1) begin            if (kd5bbe3 == 1'b1)               lsb8afd <= {yz39132{1'b0}};            else               lsb8afd <= wy15935;         end      end   end else begin      always @(*) begin         lsb8afd <= wy15935;      end   end
end
endgenerate
 shdc1a2_colorspace #(.yz39132         (yz39132       ),            .gq92cf6         (eaea539    ),            .ph329ec  (ph329ec),            .uxabeb4      (uxabeb4    ),            .yx70b70          (yx70b70        ),            .pua7b36       (pua7b36     ))     ir8a7dd (            .rstn    (rstn     ),            .clk     (clk      ),            .ce      (ngb77c       ),            .sr      (kd5bbe3       ),            .ph27078     (oh8f8b0      ),            .wwc1e36    (tj9ee2b ));
 fp81fb7_colorspace #(.yz39132         (eaea539    ),            .gq92cf6         (gq92cf6       ),            .phbf1b2      (yz39132       ),            .DOUTWIDTH      (DOUTWIDTH    ),            .sw212c2  (sw212c2),            .ph329ec  (ph329ec),            .al44ca7  (al44ca7),            .uxabeb4      (uxabeb4    ),            .ps66cfe      (ps66cfe    ),            .CPOINTS        (CPOINTS      ),            .DOUTPOINTS     (DOUTPOINTS   ),            .pua7b36       (pua7b36     ),            .nt3d9b3      (nt3d9b3    ))     ecac481 (            .rstn    (rstn     ),            .clk     (clk      ),            .ce      (ngb77c       ),            .sr      (kd5bbe3       ),            .ph27078     (bl5a3e2 ),            .wwc1e36    (wwc1e36    ));
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];wy15935<={ph27078>>1,fp2dc72[2]};bl5a3e2<={tj9ee2b>>1,fp2dc72[3]};oh8f8b0<={lsb8afd>>1,fp2dc72[4]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=ph27078[0];vk25b8e[2044]<=tj9ee2b[0];vk25b8e[2040]<=lsb8afd[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module shdc1a2_colorspace (
                 
                 clk,
                 rstn,
                 ce,
                 sr,
                 ph27078,
                 
                 wwc1e36
                 );
parameter yz39132         = 12;
parameter gq92cf6         = 12;
parameter ph329ec  = "Truncation";
parameter uxabeb4      = 3;
parameter pua7b36       = "Signed";
parameter yx70b70          = 24;
localparam  oh85b85 = (pua7b36 == "Unsigned") ? yz39132-uxabeb4 : yz39132-uxabeb4+1;
input               clk;
input               rstn;
input               ce;
input               sr;
input[yz39132-1:0]   ph27078;
output[gq92cf6-1:0]  wwc1e36;
reg                 mre20b7;
wire                ie105bc;
wire[oh85b85-1:0] nt16f08;
reg[oh85b85-1:0] ymbc23a;
reg[oh85b85-1:0] jc4d981;
reg[oh85b85-1:0] dm6cc0b;
wire[gq92cf6-1:0]    wwc1e36;
reg ngb77c;
reg kd5bbe3;
reg [yz39132 - 1 : 0] wy15935;
reg nedaaa0;
reg rgd5503;
reg [oh85b85 - 1 : 0] mr540df;
reg [oh85b85 - 1 : 0] bn37ef;
reg [oh85b85 - 1 : 0] yxc62eb;
reg [oh85b85 - 1 : 0] jr8bae8;
reg [2047:0] vk25b8e;
wire [8:0] fp2dc72;
localparam ld6e396 = 9,hb71cb6 = 32'hfdffd48b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
generate
begin   if (uxabeb4 == 0) begin         assign wwc1e36 = wy15935;   end else if (ph329ec == "Truncation") begin      assign wwc1e36 = wy15935[yz39132-1:uxabeb4];   end else begin      gbe8249_colorspace #(.yz39132  (oh85b85    ),                 .bn81692   (pua7b36    ),                 .yx70b70   (yx70b70       ))      nga8b62  (                 .rstn    (rstn    ),                 .clk     (clk     ),                 .ce      (ngb77c      ),                 .sr      (kd5bbe3      ),                 .jc4d981    (yxc62eb    ),                 .dm6cc0b    (jr8bae8    ),                 .wwc1e36    (wwc1e36    ));   end
end
endgenerate
generate
begin   if(uxabeb4 ==0 || ph329ec == "Truncation") begin      always@(*) jc4d981  <= mr540df;      always@(*) dm6cc0b  <= bn37ef;      always@(*) mre20b7  <= rgd5503;   end else begin      always @(posedge clk or negedge rstn)      begin         if (rstn == 1'b0) begin            jc4d981 <= {oh85b85{1'b0}};            dm6cc0b <= {oh85b85{1'b0}};            mre20b7  <= 1'b0;         end else if (ngb77c) begin            if (kd5bbe3) begin               jc4d981 <= {oh85b85{1'b0}};               dm6cc0b <= {oh85b85{1'b0}};               mre20b7  <= 1'b0;            end else begin               jc4d981 <= mr540df;               dm6cc0b <= bn37ef;               mre20b7  <= rgd5503;            end         end      end   end
end
endgenerate
assign ie105bc   = wy15935[yz39132-1];
generate
begin   if (pua7b36 == "Unsigned")       assign nt16f08 = {wy15935[yz39132-1:uxabeb4]};   else      assign nt16f08 = {rgd5503,wy15935[yz39132-1:uxabeb4]};
end
endgenerate
generate
begin   if (uxabeb4 > 0) begin      if (pua7b36 == "Unsigned") begin          if (ph329ec=="Rounding up") begin             always @(wy15935)               ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};         end else if (ph329ec=="Rounding away from zero") begin             always @(wy15935)               ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};         end else if (ph329ec=="Rounding towards zero") begin             always @(wy15935)            begin               if( wy15935[uxabeb4-1:0]== (1<<(uxabeb4-1)))                  ymbc23a = 0;               else                  ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};            end         end else if (ph329ec=="Convergent rounding") begin             always @(wy15935)            begin               if( wy15935[uxabeb4-1:0]== (1<<(uxabeb4-1))) begin                  if(wy15935[uxabeb4]==1)                     ymbc23a = {{(oh85b85-1){1'b0}},1'b1};                  else if(wy15935[uxabeb4]==0)                     ymbc23a = 0;               end else                  ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};            end         end      end else begin          if (ph329ec=="Rounding up") begin             always @(wy15935 or rgd5503)               ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};         end else if (ph329ec=="Rounding away from zero") begin             always @(wy15935 or rgd5503)            begin               if(rgd5503==0)                  ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};               else begin                  if( wy15935[uxabeb4-1:0]== (1<<(uxabeb4-1)))                     ymbc23a = 0;                  else                     ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};               end            end         end else if (ph329ec=="Rounding towards zero") begin             always @(wy15935 or rgd5503)            begin               if(rgd5503==0) begin                  if( wy15935[uxabeb4-1:0]== (1<<(uxabeb4-1)))                     ymbc23a = 0;                  else                     ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};               end else                  ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};            end         end else if (ph329ec=="Convergent rounding") begin             always @(wy15935 or rgd5503)            begin               if( wy15935[uxabeb4-1:0]== (1<<(uxabeb4-1))) begin                  if(wy15935[uxabeb4]==1)                     ymbc23a = {{(oh85b85-1){1'b0}},1'b1};                  else                     ymbc23a = 0;               end else                  ymbc23a = {{(oh85b85-1){1'b0}},wy15935[uxabeb4-1]};            end         end      end   end
end
endgenerate
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];wy15935<={ph27078>>1,fp2dc72[2]};nedaaa0<=fp2dc72[3];rgd5503<=fp2dc72[4];mr540df<={nt16f08>>1,fp2dc72[5]};bn37ef<={ymbc23a>>1,fp2dc72[6]};yxc62eb<={jc4d981>>1,fp2dc72[7]};jr8bae8<={dm6cc0b>>1,fp2dc72[8]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=ph27078[0];vk25b8e[2044]<=mre20b7;vk25b8e[2040]<=ie105bc;vk25b8e[2032]<=nt16f08[0];vk25b8e[2017]<=ymbc23a[0];vk25b8e[1987]<=jc4d981[0];vk25b8e[1927]<=dm6cc0b[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module fp81fb7_colorspace (
                 
                 clk,
                 rstn,
                 ce,
                 sr,
                 ph27078,
                 
                 wwc1e36
                 );
parameter yz39132         = 12;
parameter gq92cf6         = 3;
parameter phbf1b2      = 3;
parameter DOUTWIDTH      = 3;
parameter sw212c2  = 1;
parameter al44ca7  = "Saturation";
parameter ph329ec  = "Truncation";
parameter uxabeb4      = 3;
parameter ps66cfe      = 0;
parameter CPOINTS        = 0;
parameter DOUTPOINTS     = 0;
parameter pua7b36       = "Signed";
parameter nt3d9b3      = "Signed";
input                   clk;
input                   rstn;
input                   ce;
input                   sr;
input[yz39132-1:0]       ph27078;
output[DOUTWIDTH-1:0]   wwc1e36;
wire                    do4107;
wire                    zm2083a;
wire[gq92cf6-2:0]        vk20e92;
wire[gq92cf6-2:0]        ls3a495;
wire[gq92cf6-1:0]        ec9255e;
wire[gq92cf6-1:0]        wl95781;
wire[gq92cf6-1:0]        mr5e06d;
wire[gq92cf6-1:0]        hd81b60;
reg[gq92cf6-1:0]         kq6d83d;
wire[gq92cf6-1:0]        cz60f43;
reg ngb77c;
reg kd5bbe3;
reg [yz39132 - 1 : 0] wy15935;
reg tj1c9a8;
reg jce4d46;
reg [gq92cf6 - 2 : 0] ng35195;
reg [gq92cf6 - 2 : 0] me46552;
reg [gq92cf6 - 1 : 0] sj9548e;
reg [gq92cf6 - 1 : 0] tu523ae;
reg [gq92cf6 - 1 : 0] ph8eb96;
reg [gq92cf6 - 1 : 0] yzae5b5;
reg [gq92cf6 - 1 : 0] fc96d60;
reg [gq92cf6 - 1 : 0] bnb5818;
reg [2047:0] vk25b8e;
wire [12:0] fp2dc72;
localparam ld6e396 = 13,hb71cb6 = 32'hfdffe44b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
assign vk20e92  = {(gq92cf6-1){1'b1}};
assign ls3a495 = {(gq92cf6-1){1'b0}};
generate
begin   if (pua7b36 == "Unsigned") begin       if (al44ca7 == "Truncation") begin          assign hd81b60 = wy15935[gq92cf6-1:0];      end else begin          if (yz39132 == gq92cf6)            assign hd81b60 = wy15935[gq92cf6-1:0];         else begin            assign do4107 = |(wy15935[yz39132-1:gq92cf6]);            assign hd81b60 = tj1c9a8 ? {1'b1,ng35195} : wy15935[gq92cf6-1:0];         end      end   end else begin       if (nt3d9b3 == "Signed") begin         if (al44ca7=="Truncation") begin             if (uxabeb4 == 0 || ph329ec=="Truncation")               assign hd81b60 = {wy15935[yz39132-1],wy15935[gq92cf6-2:0]};            else               assign hd81b60 = {wy15935[yz39132-2],wy15935[gq92cf6-2:0]};         end else begin             if (yz39132 == gq92cf6) begin               assign hd81b60 = wy15935;            end else begin               assign do4107  = |(wy15935[yz39132-1:gq92cf6-1]);               assign zm2083a = &(wy15935[yz39132-1:gq92cf6-1]);               assign wl95781 = jce4d46 ? wy15935[gq92cf6-1:0] : {1'b1,me46552};               assign mr5e06d = tj1c9a8 ? {1'b0,ng35195} : wy15935[gq92cf6-1:0];               assign hd81b60 = wy15935[yz39132-1] ? tu523ae : ph8eb96;            end         end      end else begin          if (al44ca7 == "Truncation") begin             assign ec9255e = wy15935[gq92cf6-1:0];         end else begin             if (yz39132 == gq92cf6)               assign do4107 = 0;            else               assign do4107 = |(wy15935[yz39132-1:gq92cf6]);            assign ec9255e = tj1c9a8 ? {1'b1,ng35195} : wy15935[gq92cf6-1:0];         end         assign hd81b60 = (wy15935[yz39132-1] == 1) ? {gq92cf6{1'b0}} : sj9548e;      end   end
end
endgenerate
always @(posedge clk or negedge rstn)
begin   if (rstn == 1'b0)      kq6d83d <= {gq92cf6{1'b0}};   else if (ngb77c == 1'b1) begin      if (kd5bbe3)         kq6d83d <= {gq92cf6{1'b0}};      else         kq6d83d <= yzae5b5;   end
end
generate
begin   if (sw212c2==0) begin      assign cz60f43 = wy15935 ;   end else if(al44ca7 == "Saturation") begin      assign cz60f43 = fc96d60;   end else if((pua7b36 == "Signed") && (nt3d9b3 == "Unsigned") && (al44ca7 == "Truncation"))  begin      assign cz60f43 = fc96d60;   end else begin      assign cz60f43 = yzae5b5;   end
end
endgenerate
generate
if(DOUTPOINTS==(ps66cfe+CPOINTS)) begin   assign wwc1e36 = bnb5818;
end else if (DOUTPOINTS>(ps66cfe+CPOINTS)) begin   assign wwc1e36 = {bnb5818,{(DOUTPOINTS-(ps66cfe+CPOINTS)){1'b0}}};
end else begin   if(DOUTWIDTH<=(phbf1b2-uxabeb4))      assign wwc1e36 = bnb5818;   else begin      if (pua7b36 == "Signed")         assign wwc1e36 = {{(DOUTWIDTH-gq92cf6){bnb5818[gq92cf6-1]}},bnb5818};      else         assign wwc1e36 = {{(DOUTWIDTH-gq92cf6){1'b0}},bnb5818};   end
end
endgenerate
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];wy15935<={ph27078>>1,fp2dc72[2]};tj1c9a8<=fp2dc72[3];jce4d46<=fp2dc72[4];ng35195<={vk20e92>>1,fp2dc72[5]};me46552<={ls3a495>>1,fp2dc72[6]};sj9548e<={ec9255e>>1,fp2dc72[7]};tu523ae<={wl95781>>1,fp2dc72[8]};ph8eb96<={mr5e06d>>1,fp2dc72[9]};yzae5b5<={hd81b60>>1,fp2dc72[10]};fc96d60<={kq6d83d>>1,fp2dc72[11]};bnb5818<={cz60f43>>1,fp2dc72[12]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=ph27078[0];vk25b8e[2044]<=do4107;vk25b8e[2040]<=zm2083a;vk25b8e[2033]<=vk20e92[0];vk25b8e[2019]<=ls3a495[0];vk25b8e[1991]<=ec9255e[0];vk25b8e[1934]<=wl95781[0];vk25b8e[1821]<=mr5e06d[0];vk25b8e[1595]<=hd81b60[0];vk25b8e[1142]<=kq6d83d[0];vk25b8e[1023]<=ce;vk25b8e[237]<=cz60f43[0];end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module pf6b769_colorspace (
                     clk,   
                     rstn,
                     ce,
                     sr,
                     meef2b9,
                     din0,
                     din1,
                     din2,
                     dout0
                     );
parameter      CORETYPE          = 0;
parameter      psdaa9a        = 12;
parameter      CWIDTH            = 8;
parameter      CPOINTS           = 0;
parameter      ym3b97e      = 20;
parameter      vk2fc20    = 21;
parameter      gof081f    = 22;
parameter      DINSIGN           = "Signed";
parameter      DSPBLKMULT        = "Enable";
parameter      INSERIAL          = "Serial";
parameter      DEVICE            = "ECP2";
parameter      CV_MH             = 0;
parameter      CV_MI             = 0;
parameter      CV_MJ             = 0;
parameter      CV_MK             = 0;
parameter      CV_NH             = 0;
parameter      CV_NI             = 0;
parameter      CV_NJ             = 0;
parameter      CV_NK             = 0;
parameter      CV_PH             = 0;
parameter      CV_PI             = 0;
parameter      CV_PJ             = 0;
parameter      CV_PK             = 0;
localparam     qiadca             =  DINSIGN == "Signed" ? 1'b1 : 1'b0;
input                                     clk;
input                                     rstn;
input                                     ce;
input                                     sr;
input                                     meef2b9;
input  [psdaa9a-1:0]                   din0;
input  [psdaa9a-1:0]                   din1;
input  [psdaa9a-1:0]                   din2;
output [gof081f-1:0]               dout0;
wire   [ym3b97e-1:0]                 ld7bf5e;
wire   [ym3b97e-1:0]                 shfd7b3;
wire   [ym3b97e-1:0]                 gb5ece3;
wire   [ym3b97e-1:0]                 ecb9b35;
wire   [ym3b97e-1:0]                 zk6cd4f;
wire   [ym3b97e-1:0]                 vk353d3;
reg    [1:0]                              ksa9e9a;
reg    [CWIDTH-1:0]                       cz7a687;
reg    [CWIDTH-1:0]                       ux9a1ec;
reg    [CWIDTH-1:0]                       ou87b22;
reg    [CWIDTH-1:0]                       thec887;
reg    [CWIDTH-1:0]                       tj221f7;
reg    [CWIDTH-1:0]                       aa87df0;
reg    [ym3b97e-1:0]                 enf7c00;
reg    [ym3b97e-1:0]                 cmf0025;
reg    [ym3b97e-1:0]                 ym944;
reg    [ym3b97e-1:0]                 vk2510b;
reg    [ym3b97e-1:0]                 yma32a1;
reg    [ym3b97e-1:0]                 psca847;
reg    [ym3b97e-1:0]                 ira11d5;
reg    [vk2fc20-1:0]               qt6f1bc;
reg    [vk2fc20-1:0]               wjc6f21;
reg    [gof081f-1:0]               aabc866;
reg ngb77c;
reg kd5bbe3;
reg vka24c3;
reg [psdaa9a - 1 : 0] jc7c771;
reg [psdaa9a - 1 : 0] oh1dc57;
reg [psdaa9a - 1 : 0] jp715e2;
reg [ym3b97e - 1 : 0] kq59239;
reg [ym3b97e - 1 : 0] jc48e4c;
reg [ym3b97e - 1 : 0] ep3931b;
reg [ym3b97e - 1 : 0] ay6709c;
reg [ym3b97e - 1 : 0] blc2706;
reg [ym3b97e - 1 : 0] do9c1bf;
reg [1 : 0] ose0dfb;
reg [CWIDTH - 1 : 0] lf37ec6;
reg [CWIDTH - 1 : 0] rgfb1b7;
reg [CWIDTH - 1 : 0] enc6dde;
reg [CWIDTH - 1 : 0] lsb77a4;
reg [CWIDTH - 1 : 0] kqde91c;
reg [CWIDTH - 1 : 0] ana470b;
reg [ym3b97e - 1 : 0] rv1c2ed;
reg [ym3b97e - 1 : 0] xybb7b;
reg [ym3b97e - 1 : 0] sheded2;
reg [ym3b97e - 1 : 0] zx7b4a4;
reg [ym3b97e - 1 : 0] vk89c87;
reg [ym3b97e - 1 : 0] cm721dd;
reg [ym3b97e - 1 : 0] mg8774c;
reg [vk2fc20 - 1 : 0] irbe997;
reg [vk2fc20 - 1 : 0] swa65e3;
reg [gof081f - 1 : 0] co978c6;
reg [2047:0] vk25b8e;
wire [28:0] fp2dc72;
localparam ld6e396 = 29,hb71cb6 = 32'hfdffd14b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      ksa9e9a<= 2'b00;   end else if (ngb77c) begin      if (kd5bbe3) begin         ksa9e9a<= 2'b00;      end else if (vka24c3 ||ose0dfb==2'b10) begin         ksa9e9a<= 2'b00;      end else begin         ksa9e9a<= ose0dfb + 1'b1;      end   end
end
always @(posedge clk or negedge rstn) begin      if (!rstn) begin         cz7a687 <= {CWIDTH{1'b0}};         ou87b22 <= {CWIDTH{1'b0}};         tj221f7 <= {CWIDTH{1'b0}};         enf7c00 <= {ym3b97e{1'b0}};      end else if (ngb77c) begin         if (kd5bbe3) begin            cz7a687 <= {CWIDTH{1'b0}};            ou87b22 <= {CWIDTH{1'b0}};            tj221f7 <= {CWIDTH{1'b0}};            enf7c00 <= {ym3b97e{1'b0}};         end else begin            case (ose0dfb)               2'b00 : begin                  cz7a687 <= CV_MH;                  ou87b22 <= CV_MI;                  tj221f7 <= CV_MJ;                  enf7c00 <= CV_MK;               end               2'b01 : begin                  cz7a687 <= CV_NH;                  ou87b22 <= CV_NI;                  tj221f7 <= CV_NJ;                  enf7c00 <= CV_NK;               end               2'b10 : begin                  cz7a687 <= CV_PH;                  ou87b22 <= CV_PI;                  tj221f7 <= CV_PJ;                  enf7c00 <= CV_PK;               end               default: begin                  cz7a687 <= CV_MH;                  ou87b22 <= CV_MI;                  tj221f7 <= CV_MJ;                  enf7c00 <= CV_MK;               end            endcase         end      end
end
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      ux9a1ec  <= {CWIDTH{1'b0}};      thec887  <= {CWIDTH{1'b0}};      aa87df0  <= {CWIDTH{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         ux9a1ec  <= {CWIDTH{1'b0}};         thec887  <= {CWIDTH{1'b0}};         aa87df0  <= {CWIDTH{1'b0}};      end else begin         ux9a1ec  <= lf37ec6;         thec887  <= enc6dde;         aa87df0  <= kqde91c;      end   end
end
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      ym944 <= {ym3b97e{1'b0}};      vk2510b <= {ym3b97e{1'b0}};      cmf0025  <= {ym3b97e{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         ym944 <= {ym3b97e{1'b0}};         vk2510b <= {ym3b97e{1'b0}};         cmf0025  <= {ym3b97e{1'b0}};      end else begin         ym944 <= rv1c2ed;         vk2510b <= sheded2;         cmf0025  <= zx7b4a4;      end   end
end
generate begin   if (DSPBLKMULT == "Enable") begin         pmi_dsp_mult   #(.pmi_dataa_width           (psdaa9a     ),                          .pmi_datab_width           (CWIDTH         ),                          .pmi_additional_pipeline   (1              ),                          .pmi_input_reg             ("on"           ),                          .pmi_output_reg            ("on"           ),                          .pmi_family                (DEVICE         ),                          .pmi_gsr                   ("enable"       ),                          .pmi_source_control_a      ("parallel"     ),                          .pmi_source_control_b      ("parallel"     ),                          .pmi_reg_inputa_clk        ("CLK0"         ),                          .pmi_reg_inputa_ce         ("CE0"          ),                          .pmi_reg_inputa_rst        ("RST0"         ),                          .pmi_reg_inputb_clk        ("CLK0"         ),                          .pmi_reg_inputb_ce         ("CE0"          ),                          .pmi_reg_inputb_rst        ("RST0"         ),                          .pmi_reg_pipeline_clk      ("CLK0"         ),                          .pmi_reg_pipeline_ce       ("CE0"          ),                          .pmi_reg_pipeline_rst      ("RST0"         ),                          .pmi_reg_output_clk        ("CLK0"         ),                          .pmi_reg_output_ce         ("CE0"          ),                          .pmi_reg_output_rst        ("RST0"         ),                          .pmi_reg_signeda_clk       ("CLK0"         ),                          .pmi_reg_signeda_ce        ("CE0"          ),                          .pmi_reg_signeda_rst       ("RST0"         ),                          .pmi_reg_signedb_clk       ("CLK0"         ),                          .pmi_reg_signedb_ce        ("CE0"          ),                          .pmi_reg_signedb_rst       ("RST0"         ),                          .pmi_pipelined_mode        ("off"          ),                          .module_type               ("pmi_dsp_mult" )                         )         zx5565d  (                          .A                         (din0           ),                          .B                         (cz7a687         ),                          .SRIA                      (               ),                          .SRIB                      (               ),                          .CLK0                      (clk            ),                          .CLK1                      (clk            ),                          .CLK2                      (clk            ),                          .CLK3                      (clk            ),                          .CE0                       (ce             ),                          .CE1                       (ce             ),                          .CE2                       (ce             ),                          .CE3                       (ce             ),                          .RST0                      (~rstn          ),                          .RST1                      (~rstn          ),                          .RST2                      (~rstn          ),                          .RST3                      (~rstn          ),                          .SignA                     (qiadca          ),                          .SignB                     (1'b1           ),                          .SourceA                   (1'b0           ),                          .SourceB                   (1'b0           ),                          .P                         (ld7bf5e     ),                          .SROA                      (               ),                          .SROB                      (               ));         assign ecb9b35 = kq59239[ym3b97e-1:0];
         pmi_dsp_mult   #(.pmi_dataa_width           (psdaa9a     ),                          .pmi_datab_width           (CWIDTH         ),                          .pmi_additional_pipeline   (1              ),                          .pmi_input_reg             ("on"           ),                          .pmi_output_reg            ("on"           ),                          .pmi_family                (DEVICE         ),                          .pmi_gsr                   ("enable"       ),                          .pmi_source_control_a      ("parallel"     ),                          .pmi_source_control_b      ("parallel"     ),                          .pmi_reg_inputa_clk        ("CLK0"         ),                          .pmi_reg_inputa_ce         ("CE0"          ),                          .pmi_reg_inputa_rst        ("RST0"         ),                          .pmi_reg_inputb_clk        ("CLK0"         ),                          .pmi_reg_inputb_ce         ("CE0"          ),                          .pmi_reg_inputb_rst        ("RST0"         ),                          .pmi_reg_pipeline_clk      ("CLK0"         ),                          .pmi_reg_pipeline_ce       ("CE0"          ),                          .pmi_reg_pipeline_rst      ("RST0"         ),                          .pmi_reg_output_clk        ("CLK0"         ),                          .pmi_reg_output_ce         ("CE0"          ),                          .pmi_reg_output_rst        ("RST0"         ),                          .pmi_reg_signeda_clk       ("CLK0"         ),                          .pmi_reg_signeda_ce        ("CE0"          ),                          .pmi_reg_signeda_rst       ("RST0"         ),                          .pmi_reg_signedb_clk       ("CLK0"         ),                          .pmi_reg_signedb_ce        ("CE0"          ),                          .pmi_reg_signedb_rst       ("RST0"         ),                          .pmi_pipelined_mode        ("off"          ),                          .module_type               ("pmi_dsp_mult" )                          )         en5e7fc  (                          .A                         (din1           ),                          .B                         (ou87b22         ),                          .SRIA                      (               ),                          .SRIB                      (               ),                          .CLK0                      (clk            ),                          .CLK1                      (clk            ),                          .CLK2                      (clk            ),                          .CLK3                      (clk            ),                          .CE0                       (ce             ),                          .CE1                       (ce             ),                          .CE2                       (ce             ),                          .CE3                       (ce             ),                          .RST0                      (~rstn          ),                          .RST1                      (~rstn          ),                          .RST2                      (~rstn          ),                          .RST3                      (~rstn          ),                          .SignA                     (qiadca          ),                          .SignB                     (1'b1           ),                          .SourceA                   (1'b0           ),                          .SourceB                   (1'b0           ),                          .P                         (shfd7b3     ),                          .SROA                      (               ),                          .SROB                      (               ));         assign zk6cd4f = jc48e4c[ym3b97e-1:0];         pmi_dsp_mult   #(.pmi_dataa_width           (psdaa9a     ),                          .pmi_datab_width           (CWIDTH         ),                          .pmi_additional_pipeline   (1              ),                          .pmi_input_reg             ("on"           ),                          .pmi_output_reg            ("on"           ),                          .pmi_family                (DEVICE         ),                          .pmi_gsr                   ("enable"       ),                          .pmi_source_control_a      ("parallel"     ),                          .pmi_source_control_b      ("parallel"     ),                          .pmi_reg_inputa_clk        ("CLK0"         ),                          .pmi_reg_inputa_ce         ("CE0"          ),                          .pmi_reg_inputa_rst        ("RST0"         ),                          .pmi_reg_inputb_clk        ("CLK0"         ),                          .pmi_reg_inputb_ce         ("CE0"          ),                          .pmi_reg_inputb_rst        ("RST0"         ),                          .pmi_reg_pipeline_clk      ("CLK0"         ),                          .pmi_reg_pipeline_ce       ("CE0"          ),                          .pmi_reg_pipeline_rst      ("RST0"         ),                          .pmi_reg_output_clk        ("CLK0"         ),                          .pmi_reg_output_ce         ("CE0"          ),                          .pmi_reg_output_rst        ("RST0"         ),                          .pmi_reg_signeda_clk       ("CLK0"         ),                          .pmi_reg_signeda_ce        ("CE0"          ),                          .pmi_reg_signeda_rst       ("RST0"         ),                          .pmi_reg_signedb_clk       ("CLK0"         ),                          .pmi_reg_signedb_ce        ("CE0"          ),                          .pmi_reg_signedb_rst       ("RST0"         ),                          .pmi_pipelined_mode        ("off"          ),                          .module_type               ("pmi_dsp_mult" )                          )         gq92975  (                          .A                         (din2           ),                          .B                         (tj221f7         ),                          .SRIA                      (               ),                          .SRIB                      (               ),                          .CLK0                      (clk            ),                          .CLK1                      (clk            ),                          .CLK2                      (clk            ),                          .CLK3                      (clk            ),                          .CE0                       (ce             ),                          .CE1                       (ce             ),                          .CE2                       (ce             ),                          .CE3                       (ce             ),                          .RST0                      (~rstn          ),                          .RST1                      (~rstn          ),                          .RST2                      (~rstn          ),                          .RST3                      (~rstn          ),                          .SignA                     (qiadca          ),                          .SignB                     (1'b1           ),                          .SourceA                   (1'b0           ),                          .SourceB                   (1'b0           ),                          .P                         (gb5ece3     ),                          .SROA                      (               ),                          .SROB                      (               ));         assign vk353d3 = ep3931b[ym3b97e-1:0];   end else begin               always @(posedge clk or negedge rstn) begin                  if (!rstn) begin                     yma32a1 <= {ym3b97e{1'b0}};                     psca847 <= {ym3b97e{1'b0}};                     ira11d5 <= {ym3b97e{1'b0}};                  end else if (ngb77c) begin                     if (kd5bbe3) begin                        yma32a1 <= {ym3b97e{1'b0}};                        psca847 <= {ym3b97e{1'b0}};                        ira11d5 <= {ym3b97e{1'b0}};                     end else begin                        yma32a1 <= kq59239;                        psca847 <= jc48e4c;
                        ira11d5 <= ep3931b;                     end                  end               end                     db199ce_colorspace # (.psdaa9a                (psdaa9a          ),                              .sj39da8                 (CWIDTH              ),                              .jc76a28                     (DINSIGN             ),                              .lsa8a16                     ("Signed"            ))                    qv12a54 (.clk                       (clk                 ),                              .rstn                      (rstn                ),                              .ce                        (ngb77c                  ),                              .sr                        (kd5bbe3                  ),                              .pub26f4                  (jc7c771                ),                              .uide8d7                  (lf37ec6              ),                              .irbe63d                  (ld7bf5e          ));                     assign ecb9b35 = vk89c87[ym3b97e-1:0];                     db199ce_colorspace # (.psdaa9a                (psdaa9a          ),                              .sj39da8                 (CWIDTH              ),                              .jc76a28                     (DINSIGN             ),                              .lsa8a16                     ("Signed"            ))                    uk825f4 (.clk                       (clk                 ),                              .rstn                      (rstn                ),                              .ce                        (ngb77c                  ),                              .sr                        (kd5bbe3                  ),                              .pub26f4                  (oh1dc57                ),                              .uide8d7                  (enc6dde              ),                              .irbe63d                  (shfd7b3          ));                     assign zk6cd4f = cm721dd[ym3b97e-1:0];                     db199ce_colorspace # (.psdaa9a                (psdaa9a          ),                              .sj39da8                 (CWIDTH              ),                              .jc76a28                     (DINSIGN             ),                              .lsa8a16                     ("Signed"            ))                    vvf9c5d (.clk                       (clk                 ),                              .rstn                      (rstn                ),                              .ce                        (ngb77c                  ),                              .sr                        (kd5bbe3                  ),                              .pub26f4                  (jp715e2                ),                              .uide8d7                  (kqde91c              ),                              .irbe63d                  (gb5ece3          ));                     assign vk353d3 = mg8774c[ym3b97e-1:0];   end
end
endgenerate
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      qt6f1bc <= {vk2fc20{1'b0}};      wjc6f21 <= {vk2fc20{1'b0}};      aabc866 <= {gof081f{1'b0}};   end else if (ngb77c) begin      if (kd5bbe3) begin         qt6f1bc <= {vk2fc20{1'b0}};         wjc6f21 <= {vk2fc20{1'b0}};         aabc866 <= {gof081f{1'b0}};      end else begin         qt6f1bc <= {ay6709c[ym3b97e-1],ay6709c} + {blc2706[ym3b97e-1],blc2706};         wjc6f21 <= {do9c1bf[ym3b97e-1],do9c1bf} + {xybb7b[ym3b97e-1],xybb7b};         aabc866 <= {irbe997[vk2fc20-1],irbe997} + {swa65e3[vk2fc20-1],swa65e3};      end   end
end
assign dout0 = co978c6;
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];vka24c3<=fp2dc72[2];jc7c771<={din0>>1,fp2dc72[3]};oh1dc57<={din1>>1,fp2dc72[4]};jp715e2<={din2>>1,fp2dc72[5]};kq59239<={ld7bf5e>>1,fp2dc72[6]};jc48e4c<={shfd7b3>>1,fp2dc72[7]};ep3931b<={gb5ece3>>1,fp2dc72[8]};ay6709c<={ecb9b35>>1,fp2dc72[9]};blc2706<={zk6cd4f>>1,fp2dc72[10]};do9c1bf<={vk353d3>>1,fp2dc72[11]};ose0dfb<={ksa9e9a>>1,fp2dc72[12]};lf37ec6<={cz7a687>>1,fp2dc72[13]};rgfb1b7<={ux9a1ec>>1,fp2dc72[14]};enc6dde<={ou87b22>>1,fp2dc72[15]};lsb77a4<={thec887>>1,fp2dc72[16]};kqde91c<={tj221f7>>1,fp2dc72[17]};ana470b<={aa87df0>>1,fp2dc72[18]};rv1c2ed<={enf7c00>>1,fp2dc72[19]};xybb7b<={cmf0025>>1,fp2dc72[20]};sheded2<={ym944>>1,fp2dc72[21]};zx7b4a4<={vk2510b>>1,fp2dc72[22]};vk89c87<={yma32a1>>1,fp2dc72[23]};cm721dd<={psca847>>1,fp2dc72[24]};mg8774c<={ira11d5>>1,fp2dc72[25]};irbe997<={qt6f1bc>>1,fp2dc72[26]};swa65e3<={wjc6f21>>1,fp2dc72[27]};co978c6<={aabc866>>1,fp2dc72[28]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=meef2b9;vk25b8e[2044]<=din0[0];vk25b8e[2040]<=din1[0];vk25b8e[2033]<=din2[0];vk25b8e[2019]<=ld7bf5e[0];vk25b8e[1990]<=shfd7b3[0];vk25b8e[1981]<=wjc6f21[0];vk25b8e[1939]<=aa87df0[0];vk25b8e[1933]<=gb5ece3[0];vk25b8e[1914]<=aabc866[0];vk25b8e[1831]<=enf7c00[0];vk25b8e[1819]<=ecb9b35[0];vk25b8e[1778]<=ou87b22[0];vk25b8e[1615]<=cmf0025[0];vk25b8e[1591]<=zk6cd4f[0];vk25b8e[1508]<=thec887[0];vk25b8e[1271]<=psca847[0];vk25b8e[1182]<=ym944[0];vk25b8e[1135]<=vk353d3[0];vk25b8e[1023]<=ce;vk25b8e[990]<=qt6f1bc[0];vk25b8e[969]<=tj221f7[0];vk25b8e[889]<=ux9a1ec[0];vk25b8e[635]<=yma32a1[0];vk25b8e[495]<=ira11d5[0];vk25b8e[444]<=cz7a687[0];vk25b8e[317]<=vk2510b[0];vk25b8e[222]<=ksa9e9a[0];end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module db199ce_colorspace (
               clk,                 
               rstn,                
               ce,                  
               sr,                  
               pub26f4,            
               uide8d7,            
               
               irbe63d             
               ) ;
parameter   psdaa9a           = 8;
parameter   sj39da8            = 12;
parameter   jc76a28                = "Signed";
parameter   lsa8a16                = "Signed";
localparam  ld740ab         = psdaa9a + sj39da8 ;
input                                     clk;
input                                     rstn;
input                                     ce;
input                                     sr;
input  [psdaa9a-1:0]                   pub26f4;
input  [sj39da8-1:0]                    uide8d7;
output [ld740ab-1:0]                 irbe63d;
wire   [ld740ab-1:0]                 nt22f98 ;
reg    [psdaa9a-1:0]                   kq43b0b;
reg    [sj39da8-1:0]                    vvec2c4;
reg    [ld740ab-1:0]                 irbe63d;
reg ngb77c;
reg kd5bbe3;
reg [psdaa9a - 1 : 0] ba3f68f;
reg [sj39da8 - 1 : 0] xwda3db;
reg [ld740ab - 1 : 0] sj8f6d0;
reg [psdaa9a - 1 : 0] ykdb42f;
reg [sj39da8 - 1 : 0] psd0bc2;
reg [2047:0] vk25b8e;
wire [6:0] fp2dc72;
localparam ld6e396 = 7,hb71cb6 = 32'hfdffd48b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
      
         always @(posedge clk or negedge rstn) begin      if (!rstn) begin         kq43b0b <= {psdaa9a{1'b0}};         vvec2c4 <= {sj39da8{1'b0}};      end else if (ngb77c) begin         if (kd5bbe3) begin            kq43b0b <= {psdaa9a{1'b0}};            vvec2c4 <= {sj39da8{1'b0}};         end else begin            kq43b0b <= ba3f68f;            vvec2c4 <= xwda3db;         end      end   end   always @(posedge clk or negedge rstn) begin      if (!rstn) begin         irbe63d <= {ld740ab{1'b0}};      end else if (ngb77c) begin         if (kd5bbe3) begin            irbe63d <= {ld740ab{1'b0}};         end else begin            irbe63d <= sj8f6d0;         end      end   end
   generate begin      if (jc76a28 == "Unsigned" && lsa8a16 == "Unsigned") begin         assign nt22f98  = {{(ld740ab-psdaa9a){1'b0}},ykdb42f} * {{(ld740ab-sj39da8){1'b0}},psd0bc2};      end else if (jc76a28 == "Unsigned" && lsa8a16 == "Signed") begin         assign nt22f98  = {{(ld740ab-psdaa9a){1'b0}},ykdb42f} * {{(ld740ab-sj39da8){psd0bc2[sj39da8-1]}},psd0bc2};      end else if (jc76a28 == "Signed" && lsa8a16 == "Unsigned") begin         assign nt22f98  = {{(ld740ab-psdaa9a){ykdb42f[psdaa9a-1]}},ykdb42f} * {{(ld740ab-sj39da8){1'b0}},psd0bc2};      end else begin         assign nt22f98  = {{(ld740ab-psdaa9a){ykdb42f[psdaa9a-1]}},ykdb42f} * {{(ld740ab-sj39da8){psd0bc2[sj39da8-1]}},psd0bc2};      end   end   endgenerate
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];ba3f68f<={pub26f4>>1,fp2dc72[2]};xwda3db<={uide8d7>>1,fp2dc72[3]};sj8f6d0<={nt22f98>>1,fp2dc72[4]};ykdb42f<={kq43b0b>>1,fp2dc72[5]};psd0bc2<={vvec2c4>>1,fp2dc72[6]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=pub26f4[0];vk25b8e[2044]<=uide8d7[0];vk25b8e[2040]<=nt22f98[0];vk25b8e[2032]<=kq43b0b[0];vk25b8e[2017]<=vvec2c4[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
module su78d89_colorspace (
               
               clk,                 
               rstn,                
               ce,                  
               sr,                  
               ww4ca1b,                
               ph27078,                 
               
               dout2,               
               dout1,               
               dout0                
               );
parameter psdaa9a           = 8;
input                                     clk;
input                                     rstn;
input                                     ce;
input                                     sr;
input                                     ww4ca1b;
input  [psdaa9a-1:0]                   ph27078;
output [psdaa9a-1:0]                   dout0;
output [psdaa9a-1:0]                   dout1;
output [psdaa9a-1:0]                   dout2;
reg    [psdaa9a-1:0]                   uv65e6c;
reg    [psdaa9a-1:0]                   ho79b22;
wire   [psdaa9a-1:0]                   jc6c89f;
reg    [psdaa9a-1:0]                   dout0;
reg    [psdaa9a-1:0]                   dout1;
reg    [psdaa9a-1:0]                   dout2;
reg ngb77c;
reg kd5bbe3;
reg swbc1e4;
reg [psdaa9a - 1 : 0] wy15935;
reg [psdaa9a - 1 : 0] hoe4025;
reg [psdaa9a - 1 : 0] mg95b;
reg [psdaa9a - 1 : 0] hq256cb;
reg [2047:0] vk25b8e;
wire [6:0] fp2dc72;
localparam ld6e396 = 7,hb71cb6 = 32'hfdffd30b;
localparam [31:0] jr8e5b7 = hb71cb6;
localparam pu96df8 = hb71cb6 & 4'hf;
localparam [11:0] pub7e18 = 'h7ff;
wire [(1 << pu96df8) -1:0] off8617;
reg [ld6e396-1:0] yz185e5;
reg [pu96df8-1:0] an1796e [0:1];
reg [pu96df8-1:0] yke5ba9;
reg db2dd48;
integer vv6ea46;
integer mr75237;
assign jc6c89f = wy15935;
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      uv65e6c <= 0;      ho79b22 <= 0;   end   else if (ngb77c) begin      if (kd5bbe3) begin         uv65e6c <= 0;         ho79b22 <= 0;      end      else begin         uv65e6c <= mg95b;         ho79b22 <= hq256cb;      end   end
end
always @(posedge clk or negedge rstn) begin   if (!rstn) begin      dout0 <= 0;      dout1 <= 0;      dout2 <= 0;   end   else if (ngb77c) begin      if (kd5bbe3) begin         dout0 <= 0;         dout1 <= 0;         dout2 <= 0;      end      else if (swbc1e4) begin         dout0 <= hoe4025;         dout1 <= mg95b;         dout2 <= hq256cb;      end   end
end
always@* begin ngb77c<=fp2dc72[0];kd5bbe3<=fp2dc72[1];swbc1e4<=fp2dc72[2];wy15935<={ph27078>>1,fp2dc72[3]};hoe4025<={uv65e6c>>1,fp2dc72[4]};mg95b<={ho79b22>>1,fp2dc72[5]};hq256cb<={jc6c89f>>1,fp2dc72[6]};end
always@* begin vk25b8e[2047]<=sr;vk25b8e[2046]<=ww4ca1b;vk25b8e[2044]<=ph27078[0];vk25b8e[2040]<=uv65e6c[0];vk25b8e[2032]<=ho79b22[0];vk25b8e[2016]<=jc6c89f[0];vk25b8e[1023]<=ce;end         assign off8617 = vk25b8e,fp2dc72 = yz185e5; initial begin vv6ea46 = $fopen(".fred"); $fdisplay( vv6ea46, "%3h\n%3h", (jr8e5b7 >> 4) & pub7e18, (jr8e5b7 >> (pu96df8+4)) & pub7e18 ); $fclose(vv6ea46); $readmemh(".fred", an1796e); end always @ (off8617) begin yke5ba9 = an1796e[1]; for (mr75237=0; mr75237<ld6e396; mr75237=mr75237+1) begin yz185e5[mr75237] = off8617[yke5ba9]; db2dd48 = ^(yke5ba9 & an1796e[0]); yke5ba9 = {yke5ba9, db2dd48}; end end 
endmodule
