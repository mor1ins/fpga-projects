//////////////////////////////////////////////////////////////////////////////////
// Module Name:    i2c_ctrl 
// Description:    
// generate the instruction to config the  tvp5154/saa7129 devices iva I2C
// 0.1 --- December 18 2009 --- File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
module hdmi_i2c_ctrl (
   input  wire       rst_n      ,
   input  wire       clk        ,
   output wire       config_done,
   output reg        cmd        ,
   output reg  [6:0] addr_dev   ,
   output reg  [7:0] addr_reg_H ,
   output reg  [7:0] addr_reg_L ,
   output reg  [7:0] data_wr_H  ,
   output reg  [7:0] data_wr_L  ,
   input  wire       data_rdy   ,
   input  wire [7:0] data_rd    ,
   input  wire       i2c_done   ,
   output reg        i2c_rqt

   )/* synthesis syn_preserve=1 */
   /* synthesis syn_hier = "hard" */;


   reg               i2c_done_s1;
   reg [11:0]         step_cnt;
   wire              i2c_done_neg;

   
   parameter  
      WRITE= 1,
      READ = 0;

   
   parameter ADDR_SENSOR  =7'h3B;




   always@(posedge clk ) i2c_done_s1<=i2c_done;
   assign i2c_done_neg = !i2c_done && i2c_done_s1;
  
   always@(posedge clk or  negedge rst_n) begin
      if(!rst_n) begin
         i2c_rqt <= 0;
         step_cnt<=0;   
      end
      else if ( step_cnt<=30) begin // TBD: how many registers need to be configured.
        if(i2c_done_neg) begin
           step_cnt<=step_cnt+1; 
           i2c_rqt <= 1'b0;
        end
        else 
           i2c_rqt <= 1'b1;
      end   
      else if (i2c_done_neg)
         i2c_rqt <= 1'b0;    
   end
   
assign config_done = (step_cnt==31);
   
   always@(*) begin
         case( step_cnt)			 

 			 0:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'hC7; data_wr_H=8'h00; end // HDMI configuration
				 
			 2:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h1E; data_wr_H=8'h00; end // Power Up Transmitter
			 3:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h08; data_wr_H=8'h60; end // Input Bus/Pixel Repetition (default)
				 
			 4:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h00; data_wr_H=8'h02; end // Pixel Clock
			 5:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h01; data_wr_H=8'h3A; end // 
				 
			 6:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h02; data_wr_H=8'h70; end // Frame Rate * 100
			 7:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h03; data_wr_H=8'h17; end //

			 8:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h04; data_wr_H=8'h98; end // Pixels
			 9:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h05; data_wr_H=8'h08; end // 
				 
			 10:  begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h06; data_wr_H=8'h65; end // Lines
			 11:  begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h07; data_wr_H=8'h04; end // 	
				 
             30:   begin cmd=WRITE; addr_dev=ADDR_SENSOR; addr_reg_H=8'h1A; data_wr_H=8'h00; end
		     
            default:  begin ;end    
         endcase                                                                                            

                                                                                                            
   end                                                                                                      
                                                                                                            
                                                                                                            
endmodule                                                                                                   
                                                                                                            





















































































































































































































































































































































            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            
            