//------------------------------------------------
// USERNAME module instantiation template
//------------------------------------------------
colorspace u1_colorspace (
               .clk(clk),
               .din0(din0),
               .din1(din1),
               .din2(din2),
               .dout0(dout0),
               .dout1(dout1),
               .dout2(dout2),
               .rstn(rstn)
);
